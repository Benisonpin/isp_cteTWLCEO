magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< nwell >>
rect -1352 -1219 1352 1219
<< pmos >>
rect -1156 -1000 -1056 1000
rect -998 -1000 -898 1000
rect -840 -1000 -740 1000
rect -682 -1000 -582 1000
rect -524 -1000 -424 1000
rect -366 -1000 -266 1000
rect -208 -1000 -108 1000
rect -50 -1000 50 1000
rect 108 -1000 208 1000
rect 266 -1000 366 1000
rect 424 -1000 524 1000
rect 582 -1000 682 1000
rect 740 -1000 840 1000
rect 898 -1000 998 1000
rect 1056 -1000 1156 1000
<< pdiff >>
rect -1214 969 -1156 1000
rect -1214 935 -1202 969
rect -1168 935 -1156 969
rect -1214 901 -1156 935
rect -1214 867 -1202 901
rect -1168 867 -1156 901
rect -1214 833 -1156 867
rect -1214 799 -1202 833
rect -1168 799 -1156 833
rect -1214 765 -1156 799
rect -1214 731 -1202 765
rect -1168 731 -1156 765
rect -1214 697 -1156 731
rect -1214 663 -1202 697
rect -1168 663 -1156 697
rect -1214 629 -1156 663
rect -1214 595 -1202 629
rect -1168 595 -1156 629
rect -1214 561 -1156 595
rect -1214 527 -1202 561
rect -1168 527 -1156 561
rect -1214 493 -1156 527
rect -1214 459 -1202 493
rect -1168 459 -1156 493
rect -1214 425 -1156 459
rect -1214 391 -1202 425
rect -1168 391 -1156 425
rect -1214 357 -1156 391
rect -1214 323 -1202 357
rect -1168 323 -1156 357
rect -1214 289 -1156 323
rect -1214 255 -1202 289
rect -1168 255 -1156 289
rect -1214 221 -1156 255
rect -1214 187 -1202 221
rect -1168 187 -1156 221
rect -1214 153 -1156 187
rect -1214 119 -1202 153
rect -1168 119 -1156 153
rect -1214 85 -1156 119
rect -1214 51 -1202 85
rect -1168 51 -1156 85
rect -1214 17 -1156 51
rect -1214 -17 -1202 17
rect -1168 -17 -1156 17
rect -1214 -51 -1156 -17
rect -1214 -85 -1202 -51
rect -1168 -85 -1156 -51
rect -1214 -119 -1156 -85
rect -1214 -153 -1202 -119
rect -1168 -153 -1156 -119
rect -1214 -187 -1156 -153
rect -1214 -221 -1202 -187
rect -1168 -221 -1156 -187
rect -1214 -255 -1156 -221
rect -1214 -289 -1202 -255
rect -1168 -289 -1156 -255
rect -1214 -323 -1156 -289
rect -1214 -357 -1202 -323
rect -1168 -357 -1156 -323
rect -1214 -391 -1156 -357
rect -1214 -425 -1202 -391
rect -1168 -425 -1156 -391
rect -1214 -459 -1156 -425
rect -1214 -493 -1202 -459
rect -1168 -493 -1156 -459
rect -1214 -527 -1156 -493
rect -1214 -561 -1202 -527
rect -1168 -561 -1156 -527
rect -1214 -595 -1156 -561
rect -1214 -629 -1202 -595
rect -1168 -629 -1156 -595
rect -1214 -663 -1156 -629
rect -1214 -697 -1202 -663
rect -1168 -697 -1156 -663
rect -1214 -731 -1156 -697
rect -1214 -765 -1202 -731
rect -1168 -765 -1156 -731
rect -1214 -799 -1156 -765
rect -1214 -833 -1202 -799
rect -1168 -833 -1156 -799
rect -1214 -867 -1156 -833
rect -1214 -901 -1202 -867
rect -1168 -901 -1156 -867
rect -1214 -935 -1156 -901
rect -1214 -969 -1202 -935
rect -1168 -969 -1156 -935
rect -1214 -1000 -1156 -969
rect -1056 969 -998 1000
rect -1056 935 -1044 969
rect -1010 935 -998 969
rect -1056 901 -998 935
rect -1056 867 -1044 901
rect -1010 867 -998 901
rect -1056 833 -998 867
rect -1056 799 -1044 833
rect -1010 799 -998 833
rect -1056 765 -998 799
rect -1056 731 -1044 765
rect -1010 731 -998 765
rect -1056 697 -998 731
rect -1056 663 -1044 697
rect -1010 663 -998 697
rect -1056 629 -998 663
rect -1056 595 -1044 629
rect -1010 595 -998 629
rect -1056 561 -998 595
rect -1056 527 -1044 561
rect -1010 527 -998 561
rect -1056 493 -998 527
rect -1056 459 -1044 493
rect -1010 459 -998 493
rect -1056 425 -998 459
rect -1056 391 -1044 425
rect -1010 391 -998 425
rect -1056 357 -998 391
rect -1056 323 -1044 357
rect -1010 323 -998 357
rect -1056 289 -998 323
rect -1056 255 -1044 289
rect -1010 255 -998 289
rect -1056 221 -998 255
rect -1056 187 -1044 221
rect -1010 187 -998 221
rect -1056 153 -998 187
rect -1056 119 -1044 153
rect -1010 119 -998 153
rect -1056 85 -998 119
rect -1056 51 -1044 85
rect -1010 51 -998 85
rect -1056 17 -998 51
rect -1056 -17 -1044 17
rect -1010 -17 -998 17
rect -1056 -51 -998 -17
rect -1056 -85 -1044 -51
rect -1010 -85 -998 -51
rect -1056 -119 -998 -85
rect -1056 -153 -1044 -119
rect -1010 -153 -998 -119
rect -1056 -187 -998 -153
rect -1056 -221 -1044 -187
rect -1010 -221 -998 -187
rect -1056 -255 -998 -221
rect -1056 -289 -1044 -255
rect -1010 -289 -998 -255
rect -1056 -323 -998 -289
rect -1056 -357 -1044 -323
rect -1010 -357 -998 -323
rect -1056 -391 -998 -357
rect -1056 -425 -1044 -391
rect -1010 -425 -998 -391
rect -1056 -459 -998 -425
rect -1056 -493 -1044 -459
rect -1010 -493 -998 -459
rect -1056 -527 -998 -493
rect -1056 -561 -1044 -527
rect -1010 -561 -998 -527
rect -1056 -595 -998 -561
rect -1056 -629 -1044 -595
rect -1010 -629 -998 -595
rect -1056 -663 -998 -629
rect -1056 -697 -1044 -663
rect -1010 -697 -998 -663
rect -1056 -731 -998 -697
rect -1056 -765 -1044 -731
rect -1010 -765 -998 -731
rect -1056 -799 -998 -765
rect -1056 -833 -1044 -799
rect -1010 -833 -998 -799
rect -1056 -867 -998 -833
rect -1056 -901 -1044 -867
rect -1010 -901 -998 -867
rect -1056 -935 -998 -901
rect -1056 -969 -1044 -935
rect -1010 -969 -998 -935
rect -1056 -1000 -998 -969
rect -898 969 -840 1000
rect -898 935 -886 969
rect -852 935 -840 969
rect -898 901 -840 935
rect -898 867 -886 901
rect -852 867 -840 901
rect -898 833 -840 867
rect -898 799 -886 833
rect -852 799 -840 833
rect -898 765 -840 799
rect -898 731 -886 765
rect -852 731 -840 765
rect -898 697 -840 731
rect -898 663 -886 697
rect -852 663 -840 697
rect -898 629 -840 663
rect -898 595 -886 629
rect -852 595 -840 629
rect -898 561 -840 595
rect -898 527 -886 561
rect -852 527 -840 561
rect -898 493 -840 527
rect -898 459 -886 493
rect -852 459 -840 493
rect -898 425 -840 459
rect -898 391 -886 425
rect -852 391 -840 425
rect -898 357 -840 391
rect -898 323 -886 357
rect -852 323 -840 357
rect -898 289 -840 323
rect -898 255 -886 289
rect -852 255 -840 289
rect -898 221 -840 255
rect -898 187 -886 221
rect -852 187 -840 221
rect -898 153 -840 187
rect -898 119 -886 153
rect -852 119 -840 153
rect -898 85 -840 119
rect -898 51 -886 85
rect -852 51 -840 85
rect -898 17 -840 51
rect -898 -17 -886 17
rect -852 -17 -840 17
rect -898 -51 -840 -17
rect -898 -85 -886 -51
rect -852 -85 -840 -51
rect -898 -119 -840 -85
rect -898 -153 -886 -119
rect -852 -153 -840 -119
rect -898 -187 -840 -153
rect -898 -221 -886 -187
rect -852 -221 -840 -187
rect -898 -255 -840 -221
rect -898 -289 -886 -255
rect -852 -289 -840 -255
rect -898 -323 -840 -289
rect -898 -357 -886 -323
rect -852 -357 -840 -323
rect -898 -391 -840 -357
rect -898 -425 -886 -391
rect -852 -425 -840 -391
rect -898 -459 -840 -425
rect -898 -493 -886 -459
rect -852 -493 -840 -459
rect -898 -527 -840 -493
rect -898 -561 -886 -527
rect -852 -561 -840 -527
rect -898 -595 -840 -561
rect -898 -629 -886 -595
rect -852 -629 -840 -595
rect -898 -663 -840 -629
rect -898 -697 -886 -663
rect -852 -697 -840 -663
rect -898 -731 -840 -697
rect -898 -765 -886 -731
rect -852 -765 -840 -731
rect -898 -799 -840 -765
rect -898 -833 -886 -799
rect -852 -833 -840 -799
rect -898 -867 -840 -833
rect -898 -901 -886 -867
rect -852 -901 -840 -867
rect -898 -935 -840 -901
rect -898 -969 -886 -935
rect -852 -969 -840 -935
rect -898 -1000 -840 -969
rect -740 969 -682 1000
rect -740 935 -728 969
rect -694 935 -682 969
rect -740 901 -682 935
rect -740 867 -728 901
rect -694 867 -682 901
rect -740 833 -682 867
rect -740 799 -728 833
rect -694 799 -682 833
rect -740 765 -682 799
rect -740 731 -728 765
rect -694 731 -682 765
rect -740 697 -682 731
rect -740 663 -728 697
rect -694 663 -682 697
rect -740 629 -682 663
rect -740 595 -728 629
rect -694 595 -682 629
rect -740 561 -682 595
rect -740 527 -728 561
rect -694 527 -682 561
rect -740 493 -682 527
rect -740 459 -728 493
rect -694 459 -682 493
rect -740 425 -682 459
rect -740 391 -728 425
rect -694 391 -682 425
rect -740 357 -682 391
rect -740 323 -728 357
rect -694 323 -682 357
rect -740 289 -682 323
rect -740 255 -728 289
rect -694 255 -682 289
rect -740 221 -682 255
rect -740 187 -728 221
rect -694 187 -682 221
rect -740 153 -682 187
rect -740 119 -728 153
rect -694 119 -682 153
rect -740 85 -682 119
rect -740 51 -728 85
rect -694 51 -682 85
rect -740 17 -682 51
rect -740 -17 -728 17
rect -694 -17 -682 17
rect -740 -51 -682 -17
rect -740 -85 -728 -51
rect -694 -85 -682 -51
rect -740 -119 -682 -85
rect -740 -153 -728 -119
rect -694 -153 -682 -119
rect -740 -187 -682 -153
rect -740 -221 -728 -187
rect -694 -221 -682 -187
rect -740 -255 -682 -221
rect -740 -289 -728 -255
rect -694 -289 -682 -255
rect -740 -323 -682 -289
rect -740 -357 -728 -323
rect -694 -357 -682 -323
rect -740 -391 -682 -357
rect -740 -425 -728 -391
rect -694 -425 -682 -391
rect -740 -459 -682 -425
rect -740 -493 -728 -459
rect -694 -493 -682 -459
rect -740 -527 -682 -493
rect -740 -561 -728 -527
rect -694 -561 -682 -527
rect -740 -595 -682 -561
rect -740 -629 -728 -595
rect -694 -629 -682 -595
rect -740 -663 -682 -629
rect -740 -697 -728 -663
rect -694 -697 -682 -663
rect -740 -731 -682 -697
rect -740 -765 -728 -731
rect -694 -765 -682 -731
rect -740 -799 -682 -765
rect -740 -833 -728 -799
rect -694 -833 -682 -799
rect -740 -867 -682 -833
rect -740 -901 -728 -867
rect -694 -901 -682 -867
rect -740 -935 -682 -901
rect -740 -969 -728 -935
rect -694 -969 -682 -935
rect -740 -1000 -682 -969
rect -582 969 -524 1000
rect -582 935 -570 969
rect -536 935 -524 969
rect -582 901 -524 935
rect -582 867 -570 901
rect -536 867 -524 901
rect -582 833 -524 867
rect -582 799 -570 833
rect -536 799 -524 833
rect -582 765 -524 799
rect -582 731 -570 765
rect -536 731 -524 765
rect -582 697 -524 731
rect -582 663 -570 697
rect -536 663 -524 697
rect -582 629 -524 663
rect -582 595 -570 629
rect -536 595 -524 629
rect -582 561 -524 595
rect -582 527 -570 561
rect -536 527 -524 561
rect -582 493 -524 527
rect -582 459 -570 493
rect -536 459 -524 493
rect -582 425 -524 459
rect -582 391 -570 425
rect -536 391 -524 425
rect -582 357 -524 391
rect -582 323 -570 357
rect -536 323 -524 357
rect -582 289 -524 323
rect -582 255 -570 289
rect -536 255 -524 289
rect -582 221 -524 255
rect -582 187 -570 221
rect -536 187 -524 221
rect -582 153 -524 187
rect -582 119 -570 153
rect -536 119 -524 153
rect -582 85 -524 119
rect -582 51 -570 85
rect -536 51 -524 85
rect -582 17 -524 51
rect -582 -17 -570 17
rect -536 -17 -524 17
rect -582 -51 -524 -17
rect -582 -85 -570 -51
rect -536 -85 -524 -51
rect -582 -119 -524 -85
rect -582 -153 -570 -119
rect -536 -153 -524 -119
rect -582 -187 -524 -153
rect -582 -221 -570 -187
rect -536 -221 -524 -187
rect -582 -255 -524 -221
rect -582 -289 -570 -255
rect -536 -289 -524 -255
rect -582 -323 -524 -289
rect -582 -357 -570 -323
rect -536 -357 -524 -323
rect -582 -391 -524 -357
rect -582 -425 -570 -391
rect -536 -425 -524 -391
rect -582 -459 -524 -425
rect -582 -493 -570 -459
rect -536 -493 -524 -459
rect -582 -527 -524 -493
rect -582 -561 -570 -527
rect -536 -561 -524 -527
rect -582 -595 -524 -561
rect -582 -629 -570 -595
rect -536 -629 -524 -595
rect -582 -663 -524 -629
rect -582 -697 -570 -663
rect -536 -697 -524 -663
rect -582 -731 -524 -697
rect -582 -765 -570 -731
rect -536 -765 -524 -731
rect -582 -799 -524 -765
rect -582 -833 -570 -799
rect -536 -833 -524 -799
rect -582 -867 -524 -833
rect -582 -901 -570 -867
rect -536 -901 -524 -867
rect -582 -935 -524 -901
rect -582 -969 -570 -935
rect -536 -969 -524 -935
rect -582 -1000 -524 -969
rect -424 969 -366 1000
rect -424 935 -412 969
rect -378 935 -366 969
rect -424 901 -366 935
rect -424 867 -412 901
rect -378 867 -366 901
rect -424 833 -366 867
rect -424 799 -412 833
rect -378 799 -366 833
rect -424 765 -366 799
rect -424 731 -412 765
rect -378 731 -366 765
rect -424 697 -366 731
rect -424 663 -412 697
rect -378 663 -366 697
rect -424 629 -366 663
rect -424 595 -412 629
rect -378 595 -366 629
rect -424 561 -366 595
rect -424 527 -412 561
rect -378 527 -366 561
rect -424 493 -366 527
rect -424 459 -412 493
rect -378 459 -366 493
rect -424 425 -366 459
rect -424 391 -412 425
rect -378 391 -366 425
rect -424 357 -366 391
rect -424 323 -412 357
rect -378 323 -366 357
rect -424 289 -366 323
rect -424 255 -412 289
rect -378 255 -366 289
rect -424 221 -366 255
rect -424 187 -412 221
rect -378 187 -366 221
rect -424 153 -366 187
rect -424 119 -412 153
rect -378 119 -366 153
rect -424 85 -366 119
rect -424 51 -412 85
rect -378 51 -366 85
rect -424 17 -366 51
rect -424 -17 -412 17
rect -378 -17 -366 17
rect -424 -51 -366 -17
rect -424 -85 -412 -51
rect -378 -85 -366 -51
rect -424 -119 -366 -85
rect -424 -153 -412 -119
rect -378 -153 -366 -119
rect -424 -187 -366 -153
rect -424 -221 -412 -187
rect -378 -221 -366 -187
rect -424 -255 -366 -221
rect -424 -289 -412 -255
rect -378 -289 -366 -255
rect -424 -323 -366 -289
rect -424 -357 -412 -323
rect -378 -357 -366 -323
rect -424 -391 -366 -357
rect -424 -425 -412 -391
rect -378 -425 -366 -391
rect -424 -459 -366 -425
rect -424 -493 -412 -459
rect -378 -493 -366 -459
rect -424 -527 -366 -493
rect -424 -561 -412 -527
rect -378 -561 -366 -527
rect -424 -595 -366 -561
rect -424 -629 -412 -595
rect -378 -629 -366 -595
rect -424 -663 -366 -629
rect -424 -697 -412 -663
rect -378 -697 -366 -663
rect -424 -731 -366 -697
rect -424 -765 -412 -731
rect -378 -765 -366 -731
rect -424 -799 -366 -765
rect -424 -833 -412 -799
rect -378 -833 -366 -799
rect -424 -867 -366 -833
rect -424 -901 -412 -867
rect -378 -901 -366 -867
rect -424 -935 -366 -901
rect -424 -969 -412 -935
rect -378 -969 -366 -935
rect -424 -1000 -366 -969
rect -266 969 -208 1000
rect -266 935 -254 969
rect -220 935 -208 969
rect -266 901 -208 935
rect -266 867 -254 901
rect -220 867 -208 901
rect -266 833 -208 867
rect -266 799 -254 833
rect -220 799 -208 833
rect -266 765 -208 799
rect -266 731 -254 765
rect -220 731 -208 765
rect -266 697 -208 731
rect -266 663 -254 697
rect -220 663 -208 697
rect -266 629 -208 663
rect -266 595 -254 629
rect -220 595 -208 629
rect -266 561 -208 595
rect -266 527 -254 561
rect -220 527 -208 561
rect -266 493 -208 527
rect -266 459 -254 493
rect -220 459 -208 493
rect -266 425 -208 459
rect -266 391 -254 425
rect -220 391 -208 425
rect -266 357 -208 391
rect -266 323 -254 357
rect -220 323 -208 357
rect -266 289 -208 323
rect -266 255 -254 289
rect -220 255 -208 289
rect -266 221 -208 255
rect -266 187 -254 221
rect -220 187 -208 221
rect -266 153 -208 187
rect -266 119 -254 153
rect -220 119 -208 153
rect -266 85 -208 119
rect -266 51 -254 85
rect -220 51 -208 85
rect -266 17 -208 51
rect -266 -17 -254 17
rect -220 -17 -208 17
rect -266 -51 -208 -17
rect -266 -85 -254 -51
rect -220 -85 -208 -51
rect -266 -119 -208 -85
rect -266 -153 -254 -119
rect -220 -153 -208 -119
rect -266 -187 -208 -153
rect -266 -221 -254 -187
rect -220 -221 -208 -187
rect -266 -255 -208 -221
rect -266 -289 -254 -255
rect -220 -289 -208 -255
rect -266 -323 -208 -289
rect -266 -357 -254 -323
rect -220 -357 -208 -323
rect -266 -391 -208 -357
rect -266 -425 -254 -391
rect -220 -425 -208 -391
rect -266 -459 -208 -425
rect -266 -493 -254 -459
rect -220 -493 -208 -459
rect -266 -527 -208 -493
rect -266 -561 -254 -527
rect -220 -561 -208 -527
rect -266 -595 -208 -561
rect -266 -629 -254 -595
rect -220 -629 -208 -595
rect -266 -663 -208 -629
rect -266 -697 -254 -663
rect -220 -697 -208 -663
rect -266 -731 -208 -697
rect -266 -765 -254 -731
rect -220 -765 -208 -731
rect -266 -799 -208 -765
rect -266 -833 -254 -799
rect -220 -833 -208 -799
rect -266 -867 -208 -833
rect -266 -901 -254 -867
rect -220 -901 -208 -867
rect -266 -935 -208 -901
rect -266 -969 -254 -935
rect -220 -969 -208 -935
rect -266 -1000 -208 -969
rect -108 969 -50 1000
rect -108 935 -96 969
rect -62 935 -50 969
rect -108 901 -50 935
rect -108 867 -96 901
rect -62 867 -50 901
rect -108 833 -50 867
rect -108 799 -96 833
rect -62 799 -50 833
rect -108 765 -50 799
rect -108 731 -96 765
rect -62 731 -50 765
rect -108 697 -50 731
rect -108 663 -96 697
rect -62 663 -50 697
rect -108 629 -50 663
rect -108 595 -96 629
rect -62 595 -50 629
rect -108 561 -50 595
rect -108 527 -96 561
rect -62 527 -50 561
rect -108 493 -50 527
rect -108 459 -96 493
rect -62 459 -50 493
rect -108 425 -50 459
rect -108 391 -96 425
rect -62 391 -50 425
rect -108 357 -50 391
rect -108 323 -96 357
rect -62 323 -50 357
rect -108 289 -50 323
rect -108 255 -96 289
rect -62 255 -50 289
rect -108 221 -50 255
rect -108 187 -96 221
rect -62 187 -50 221
rect -108 153 -50 187
rect -108 119 -96 153
rect -62 119 -50 153
rect -108 85 -50 119
rect -108 51 -96 85
rect -62 51 -50 85
rect -108 17 -50 51
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -51 -50 -17
rect -108 -85 -96 -51
rect -62 -85 -50 -51
rect -108 -119 -50 -85
rect -108 -153 -96 -119
rect -62 -153 -50 -119
rect -108 -187 -50 -153
rect -108 -221 -96 -187
rect -62 -221 -50 -187
rect -108 -255 -50 -221
rect -108 -289 -96 -255
rect -62 -289 -50 -255
rect -108 -323 -50 -289
rect -108 -357 -96 -323
rect -62 -357 -50 -323
rect -108 -391 -50 -357
rect -108 -425 -96 -391
rect -62 -425 -50 -391
rect -108 -459 -50 -425
rect -108 -493 -96 -459
rect -62 -493 -50 -459
rect -108 -527 -50 -493
rect -108 -561 -96 -527
rect -62 -561 -50 -527
rect -108 -595 -50 -561
rect -108 -629 -96 -595
rect -62 -629 -50 -595
rect -108 -663 -50 -629
rect -108 -697 -96 -663
rect -62 -697 -50 -663
rect -108 -731 -50 -697
rect -108 -765 -96 -731
rect -62 -765 -50 -731
rect -108 -799 -50 -765
rect -108 -833 -96 -799
rect -62 -833 -50 -799
rect -108 -867 -50 -833
rect -108 -901 -96 -867
rect -62 -901 -50 -867
rect -108 -935 -50 -901
rect -108 -969 -96 -935
rect -62 -969 -50 -935
rect -108 -1000 -50 -969
rect 50 969 108 1000
rect 50 935 62 969
rect 96 935 108 969
rect 50 901 108 935
rect 50 867 62 901
rect 96 867 108 901
rect 50 833 108 867
rect 50 799 62 833
rect 96 799 108 833
rect 50 765 108 799
rect 50 731 62 765
rect 96 731 108 765
rect 50 697 108 731
rect 50 663 62 697
rect 96 663 108 697
rect 50 629 108 663
rect 50 595 62 629
rect 96 595 108 629
rect 50 561 108 595
rect 50 527 62 561
rect 96 527 108 561
rect 50 493 108 527
rect 50 459 62 493
rect 96 459 108 493
rect 50 425 108 459
rect 50 391 62 425
rect 96 391 108 425
rect 50 357 108 391
rect 50 323 62 357
rect 96 323 108 357
rect 50 289 108 323
rect 50 255 62 289
rect 96 255 108 289
rect 50 221 108 255
rect 50 187 62 221
rect 96 187 108 221
rect 50 153 108 187
rect 50 119 62 153
rect 96 119 108 153
rect 50 85 108 119
rect 50 51 62 85
rect 96 51 108 85
rect 50 17 108 51
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -51 108 -17
rect 50 -85 62 -51
rect 96 -85 108 -51
rect 50 -119 108 -85
rect 50 -153 62 -119
rect 96 -153 108 -119
rect 50 -187 108 -153
rect 50 -221 62 -187
rect 96 -221 108 -187
rect 50 -255 108 -221
rect 50 -289 62 -255
rect 96 -289 108 -255
rect 50 -323 108 -289
rect 50 -357 62 -323
rect 96 -357 108 -323
rect 50 -391 108 -357
rect 50 -425 62 -391
rect 96 -425 108 -391
rect 50 -459 108 -425
rect 50 -493 62 -459
rect 96 -493 108 -459
rect 50 -527 108 -493
rect 50 -561 62 -527
rect 96 -561 108 -527
rect 50 -595 108 -561
rect 50 -629 62 -595
rect 96 -629 108 -595
rect 50 -663 108 -629
rect 50 -697 62 -663
rect 96 -697 108 -663
rect 50 -731 108 -697
rect 50 -765 62 -731
rect 96 -765 108 -731
rect 50 -799 108 -765
rect 50 -833 62 -799
rect 96 -833 108 -799
rect 50 -867 108 -833
rect 50 -901 62 -867
rect 96 -901 108 -867
rect 50 -935 108 -901
rect 50 -969 62 -935
rect 96 -969 108 -935
rect 50 -1000 108 -969
rect 208 969 266 1000
rect 208 935 220 969
rect 254 935 266 969
rect 208 901 266 935
rect 208 867 220 901
rect 254 867 266 901
rect 208 833 266 867
rect 208 799 220 833
rect 254 799 266 833
rect 208 765 266 799
rect 208 731 220 765
rect 254 731 266 765
rect 208 697 266 731
rect 208 663 220 697
rect 254 663 266 697
rect 208 629 266 663
rect 208 595 220 629
rect 254 595 266 629
rect 208 561 266 595
rect 208 527 220 561
rect 254 527 266 561
rect 208 493 266 527
rect 208 459 220 493
rect 254 459 266 493
rect 208 425 266 459
rect 208 391 220 425
rect 254 391 266 425
rect 208 357 266 391
rect 208 323 220 357
rect 254 323 266 357
rect 208 289 266 323
rect 208 255 220 289
rect 254 255 266 289
rect 208 221 266 255
rect 208 187 220 221
rect 254 187 266 221
rect 208 153 266 187
rect 208 119 220 153
rect 254 119 266 153
rect 208 85 266 119
rect 208 51 220 85
rect 254 51 266 85
rect 208 17 266 51
rect 208 -17 220 17
rect 254 -17 266 17
rect 208 -51 266 -17
rect 208 -85 220 -51
rect 254 -85 266 -51
rect 208 -119 266 -85
rect 208 -153 220 -119
rect 254 -153 266 -119
rect 208 -187 266 -153
rect 208 -221 220 -187
rect 254 -221 266 -187
rect 208 -255 266 -221
rect 208 -289 220 -255
rect 254 -289 266 -255
rect 208 -323 266 -289
rect 208 -357 220 -323
rect 254 -357 266 -323
rect 208 -391 266 -357
rect 208 -425 220 -391
rect 254 -425 266 -391
rect 208 -459 266 -425
rect 208 -493 220 -459
rect 254 -493 266 -459
rect 208 -527 266 -493
rect 208 -561 220 -527
rect 254 -561 266 -527
rect 208 -595 266 -561
rect 208 -629 220 -595
rect 254 -629 266 -595
rect 208 -663 266 -629
rect 208 -697 220 -663
rect 254 -697 266 -663
rect 208 -731 266 -697
rect 208 -765 220 -731
rect 254 -765 266 -731
rect 208 -799 266 -765
rect 208 -833 220 -799
rect 254 -833 266 -799
rect 208 -867 266 -833
rect 208 -901 220 -867
rect 254 -901 266 -867
rect 208 -935 266 -901
rect 208 -969 220 -935
rect 254 -969 266 -935
rect 208 -1000 266 -969
rect 366 969 424 1000
rect 366 935 378 969
rect 412 935 424 969
rect 366 901 424 935
rect 366 867 378 901
rect 412 867 424 901
rect 366 833 424 867
rect 366 799 378 833
rect 412 799 424 833
rect 366 765 424 799
rect 366 731 378 765
rect 412 731 424 765
rect 366 697 424 731
rect 366 663 378 697
rect 412 663 424 697
rect 366 629 424 663
rect 366 595 378 629
rect 412 595 424 629
rect 366 561 424 595
rect 366 527 378 561
rect 412 527 424 561
rect 366 493 424 527
rect 366 459 378 493
rect 412 459 424 493
rect 366 425 424 459
rect 366 391 378 425
rect 412 391 424 425
rect 366 357 424 391
rect 366 323 378 357
rect 412 323 424 357
rect 366 289 424 323
rect 366 255 378 289
rect 412 255 424 289
rect 366 221 424 255
rect 366 187 378 221
rect 412 187 424 221
rect 366 153 424 187
rect 366 119 378 153
rect 412 119 424 153
rect 366 85 424 119
rect 366 51 378 85
rect 412 51 424 85
rect 366 17 424 51
rect 366 -17 378 17
rect 412 -17 424 17
rect 366 -51 424 -17
rect 366 -85 378 -51
rect 412 -85 424 -51
rect 366 -119 424 -85
rect 366 -153 378 -119
rect 412 -153 424 -119
rect 366 -187 424 -153
rect 366 -221 378 -187
rect 412 -221 424 -187
rect 366 -255 424 -221
rect 366 -289 378 -255
rect 412 -289 424 -255
rect 366 -323 424 -289
rect 366 -357 378 -323
rect 412 -357 424 -323
rect 366 -391 424 -357
rect 366 -425 378 -391
rect 412 -425 424 -391
rect 366 -459 424 -425
rect 366 -493 378 -459
rect 412 -493 424 -459
rect 366 -527 424 -493
rect 366 -561 378 -527
rect 412 -561 424 -527
rect 366 -595 424 -561
rect 366 -629 378 -595
rect 412 -629 424 -595
rect 366 -663 424 -629
rect 366 -697 378 -663
rect 412 -697 424 -663
rect 366 -731 424 -697
rect 366 -765 378 -731
rect 412 -765 424 -731
rect 366 -799 424 -765
rect 366 -833 378 -799
rect 412 -833 424 -799
rect 366 -867 424 -833
rect 366 -901 378 -867
rect 412 -901 424 -867
rect 366 -935 424 -901
rect 366 -969 378 -935
rect 412 -969 424 -935
rect 366 -1000 424 -969
rect 524 969 582 1000
rect 524 935 536 969
rect 570 935 582 969
rect 524 901 582 935
rect 524 867 536 901
rect 570 867 582 901
rect 524 833 582 867
rect 524 799 536 833
rect 570 799 582 833
rect 524 765 582 799
rect 524 731 536 765
rect 570 731 582 765
rect 524 697 582 731
rect 524 663 536 697
rect 570 663 582 697
rect 524 629 582 663
rect 524 595 536 629
rect 570 595 582 629
rect 524 561 582 595
rect 524 527 536 561
rect 570 527 582 561
rect 524 493 582 527
rect 524 459 536 493
rect 570 459 582 493
rect 524 425 582 459
rect 524 391 536 425
rect 570 391 582 425
rect 524 357 582 391
rect 524 323 536 357
rect 570 323 582 357
rect 524 289 582 323
rect 524 255 536 289
rect 570 255 582 289
rect 524 221 582 255
rect 524 187 536 221
rect 570 187 582 221
rect 524 153 582 187
rect 524 119 536 153
rect 570 119 582 153
rect 524 85 582 119
rect 524 51 536 85
rect 570 51 582 85
rect 524 17 582 51
rect 524 -17 536 17
rect 570 -17 582 17
rect 524 -51 582 -17
rect 524 -85 536 -51
rect 570 -85 582 -51
rect 524 -119 582 -85
rect 524 -153 536 -119
rect 570 -153 582 -119
rect 524 -187 582 -153
rect 524 -221 536 -187
rect 570 -221 582 -187
rect 524 -255 582 -221
rect 524 -289 536 -255
rect 570 -289 582 -255
rect 524 -323 582 -289
rect 524 -357 536 -323
rect 570 -357 582 -323
rect 524 -391 582 -357
rect 524 -425 536 -391
rect 570 -425 582 -391
rect 524 -459 582 -425
rect 524 -493 536 -459
rect 570 -493 582 -459
rect 524 -527 582 -493
rect 524 -561 536 -527
rect 570 -561 582 -527
rect 524 -595 582 -561
rect 524 -629 536 -595
rect 570 -629 582 -595
rect 524 -663 582 -629
rect 524 -697 536 -663
rect 570 -697 582 -663
rect 524 -731 582 -697
rect 524 -765 536 -731
rect 570 -765 582 -731
rect 524 -799 582 -765
rect 524 -833 536 -799
rect 570 -833 582 -799
rect 524 -867 582 -833
rect 524 -901 536 -867
rect 570 -901 582 -867
rect 524 -935 582 -901
rect 524 -969 536 -935
rect 570 -969 582 -935
rect 524 -1000 582 -969
rect 682 969 740 1000
rect 682 935 694 969
rect 728 935 740 969
rect 682 901 740 935
rect 682 867 694 901
rect 728 867 740 901
rect 682 833 740 867
rect 682 799 694 833
rect 728 799 740 833
rect 682 765 740 799
rect 682 731 694 765
rect 728 731 740 765
rect 682 697 740 731
rect 682 663 694 697
rect 728 663 740 697
rect 682 629 740 663
rect 682 595 694 629
rect 728 595 740 629
rect 682 561 740 595
rect 682 527 694 561
rect 728 527 740 561
rect 682 493 740 527
rect 682 459 694 493
rect 728 459 740 493
rect 682 425 740 459
rect 682 391 694 425
rect 728 391 740 425
rect 682 357 740 391
rect 682 323 694 357
rect 728 323 740 357
rect 682 289 740 323
rect 682 255 694 289
rect 728 255 740 289
rect 682 221 740 255
rect 682 187 694 221
rect 728 187 740 221
rect 682 153 740 187
rect 682 119 694 153
rect 728 119 740 153
rect 682 85 740 119
rect 682 51 694 85
rect 728 51 740 85
rect 682 17 740 51
rect 682 -17 694 17
rect 728 -17 740 17
rect 682 -51 740 -17
rect 682 -85 694 -51
rect 728 -85 740 -51
rect 682 -119 740 -85
rect 682 -153 694 -119
rect 728 -153 740 -119
rect 682 -187 740 -153
rect 682 -221 694 -187
rect 728 -221 740 -187
rect 682 -255 740 -221
rect 682 -289 694 -255
rect 728 -289 740 -255
rect 682 -323 740 -289
rect 682 -357 694 -323
rect 728 -357 740 -323
rect 682 -391 740 -357
rect 682 -425 694 -391
rect 728 -425 740 -391
rect 682 -459 740 -425
rect 682 -493 694 -459
rect 728 -493 740 -459
rect 682 -527 740 -493
rect 682 -561 694 -527
rect 728 -561 740 -527
rect 682 -595 740 -561
rect 682 -629 694 -595
rect 728 -629 740 -595
rect 682 -663 740 -629
rect 682 -697 694 -663
rect 728 -697 740 -663
rect 682 -731 740 -697
rect 682 -765 694 -731
rect 728 -765 740 -731
rect 682 -799 740 -765
rect 682 -833 694 -799
rect 728 -833 740 -799
rect 682 -867 740 -833
rect 682 -901 694 -867
rect 728 -901 740 -867
rect 682 -935 740 -901
rect 682 -969 694 -935
rect 728 -969 740 -935
rect 682 -1000 740 -969
rect 840 969 898 1000
rect 840 935 852 969
rect 886 935 898 969
rect 840 901 898 935
rect 840 867 852 901
rect 886 867 898 901
rect 840 833 898 867
rect 840 799 852 833
rect 886 799 898 833
rect 840 765 898 799
rect 840 731 852 765
rect 886 731 898 765
rect 840 697 898 731
rect 840 663 852 697
rect 886 663 898 697
rect 840 629 898 663
rect 840 595 852 629
rect 886 595 898 629
rect 840 561 898 595
rect 840 527 852 561
rect 886 527 898 561
rect 840 493 898 527
rect 840 459 852 493
rect 886 459 898 493
rect 840 425 898 459
rect 840 391 852 425
rect 886 391 898 425
rect 840 357 898 391
rect 840 323 852 357
rect 886 323 898 357
rect 840 289 898 323
rect 840 255 852 289
rect 886 255 898 289
rect 840 221 898 255
rect 840 187 852 221
rect 886 187 898 221
rect 840 153 898 187
rect 840 119 852 153
rect 886 119 898 153
rect 840 85 898 119
rect 840 51 852 85
rect 886 51 898 85
rect 840 17 898 51
rect 840 -17 852 17
rect 886 -17 898 17
rect 840 -51 898 -17
rect 840 -85 852 -51
rect 886 -85 898 -51
rect 840 -119 898 -85
rect 840 -153 852 -119
rect 886 -153 898 -119
rect 840 -187 898 -153
rect 840 -221 852 -187
rect 886 -221 898 -187
rect 840 -255 898 -221
rect 840 -289 852 -255
rect 886 -289 898 -255
rect 840 -323 898 -289
rect 840 -357 852 -323
rect 886 -357 898 -323
rect 840 -391 898 -357
rect 840 -425 852 -391
rect 886 -425 898 -391
rect 840 -459 898 -425
rect 840 -493 852 -459
rect 886 -493 898 -459
rect 840 -527 898 -493
rect 840 -561 852 -527
rect 886 -561 898 -527
rect 840 -595 898 -561
rect 840 -629 852 -595
rect 886 -629 898 -595
rect 840 -663 898 -629
rect 840 -697 852 -663
rect 886 -697 898 -663
rect 840 -731 898 -697
rect 840 -765 852 -731
rect 886 -765 898 -731
rect 840 -799 898 -765
rect 840 -833 852 -799
rect 886 -833 898 -799
rect 840 -867 898 -833
rect 840 -901 852 -867
rect 886 -901 898 -867
rect 840 -935 898 -901
rect 840 -969 852 -935
rect 886 -969 898 -935
rect 840 -1000 898 -969
rect 998 969 1056 1000
rect 998 935 1010 969
rect 1044 935 1056 969
rect 998 901 1056 935
rect 998 867 1010 901
rect 1044 867 1056 901
rect 998 833 1056 867
rect 998 799 1010 833
rect 1044 799 1056 833
rect 998 765 1056 799
rect 998 731 1010 765
rect 1044 731 1056 765
rect 998 697 1056 731
rect 998 663 1010 697
rect 1044 663 1056 697
rect 998 629 1056 663
rect 998 595 1010 629
rect 1044 595 1056 629
rect 998 561 1056 595
rect 998 527 1010 561
rect 1044 527 1056 561
rect 998 493 1056 527
rect 998 459 1010 493
rect 1044 459 1056 493
rect 998 425 1056 459
rect 998 391 1010 425
rect 1044 391 1056 425
rect 998 357 1056 391
rect 998 323 1010 357
rect 1044 323 1056 357
rect 998 289 1056 323
rect 998 255 1010 289
rect 1044 255 1056 289
rect 998 221 1056 255
rect 998 187 1010 221
rect 1044 187 1056 221
rect 998 153 1056 187
rect 998 119 1010 153
rect 1044 119 1056 153
rect 998 85 1056 119
rect 998 51 1010 85
rect 1044 51 1056 85
rect 998 17 1056 51
rect 998 -17 1010 17
rect 1044 -17 1056 17
rect 998 -51 1056 -17
rect 998 -85 1010 -51
rect 1044 -85 1056 -51
rect 998 -119 1056 -85
rect 998 -153 1010 -119
rect 1044 -153 1056 -119
rect 998 -187 1056 -153
rect 998 -221 1010 -187
rect 1044 -221 1056 -187
rect 998 -255 1056 -221
rect 998 -289 1010 -255
rect 1044 -289 1056 -255
rect 998 -323 1056 -289
rect 998 -357 1010 -323
rect 1044 -357 1056 -323
rect 998 -391 1056 -357
rect 998 -425 1010 -391
rect 1044 -425 1056 -391
rect 998 -459 1056 -425
rect 998 -493 1010 -459
rect 1044 -493 1056 -459
rect 998 -527 1056 -493
rect 998 -561 1010 -527
rect 1044 -561 1056 -527
rect 998 -595 1056 -561
rect 998 -629 1010 -595
rect 1044 -629 1056 -595
rect 998 -663 1056 -629
rect 998 -697 1010 -663
rect 1044 -697 1056 -663
rect 998 -731 1056 -697
rect 998 -765 1010 -731
rect 1044 -765 1056 -731
rect 998 -799 1056 -765
rect 998 -833 1010 -799
rect 1044 -833 1056 -799
rect 998 -867 1056 -833
rect 998 -901 1010 -867
rect 1044 -901 1056 -867
rect 998 -935 1056 -901
rect 998 -969 1010 -935
rect 1044 -969 1056 -935
rect 998 -1000 1056 -969
rect 1156 969 1214 1000
rect 1156 935 1168 969
rect 1202 935 1214 969
rect 1156 901 1214 935
rect 1156 867 1168 901
rect 1202 867 1214 901
rect 1156 833 1214 867
rect 1156 799 1168 833
rect 1202 799 1214 833
rect 1156 765 1214 799
rect 1156 731 1168 765
rect 1202 731 1214 765
rect 1156 697 1214 731
rect 1156 663 1168 697
rect 1202 663 1214 697
rect 1156 629 1214 663
rect 1156 595 1168 629
rect 1202 595 1214 629
rect 1156 561 1214 595
rect 1156 527 1168 561
rect 1202 527 1214 561
rect 1156 493 1214 527
rect 1156 459 1168 493
rect 1202 459 1214 493
rect 1156 425 1214 459
rect 1156 391 1168 425
rect 1202 391 1214 425
rect 1156 357 1214 391
rect 1156 323 1168 357
rect 1202 323 1214 357
rect 1156 289 1214 323
rect 1156 255 1168 289
rect 1202 255 1214 289
rect 1156 221 1214 255
rect 1156 187 1168 221
rect 1202 187 1214 221
rect 1156 153 1214 187
rect 1156 119 1168 153
rect 1202 119 1214 153
rect 1156 85 1214 119
rect 1156 51 1168 85
rect 1202 51 1214 85
rect 1156 17 1214 51
rect 1156 -17 1168 17
rect 1202 -17 1214 17
rect 1156 -51 1214 -17
rect 1156 -85 1168 -51
rect 1202 -85 1214 -51
rect 1156 -119 1214 -85
rect 1156 -153 1168 -119
rect 1202 -153 1214 -119
rect 1156 -187 1214 -153
rect 1156 -221 1168 -187
rect 1202 -221 1214 -187
rect 1156 -255 1214 -221
rect 1156 -289 1168 -255
rect 1202 -289 1214 -255
rect 1156 -323 1214 -289
rect 1156 -357 1168 -323
rect 1202 -357 1214 -323
rect 1156 -391 1214 -357
rect 1156 -425 1168 -391
rect 1202 -425 1214 -391
rect 1156 -459 1214 -425
rect 1156 -493 1168 -459
rect 1202 -493 1214 -459
rect 1156 -527 1214 -493
rect 1156 -561 1168 -527
rect 1202 -561 1214 -527
rect 1156 -595 1214 -561
rect 1156 -629 1168 -595
rect 1202 -629 1214 -595
rect 1156 -663 1214 -629
rect 1156 -697 1168 -663
rect 1202 -697 1214 -663
rect 1156 -731 1214 -697
rect 1156 -765 1168 -731
rect 1202 -765 1214 -731
rect 1156 -799 1214 -765
rect 1156 -833 1168 -799
rect 1202 -833 1214 -799
rect 1156 -867 1214 -833
rect 1156 -901 1168 -867
rect 1202 -901 1214 -867
rect 1156 -935 1214 -901
rect 1156 -969 1168 -935
rect 1202 -969 1214 -935
rect 1156 -1000 1214 -969
<< pdiffc >>
rect -1202 935 -1168 969
rect -1202 867 -1168 901
rect -1202 799 -1168 833
rect -1202 731 -1168 765
rect -1202 663 -1168 697
rect -1202 595 -1168 629
rect -1202 527 -1168 561
rect -1202 459 -1168 493
rect -1202 391 -1168 425
rect -1202 323 -1168 357
rect -1202 255 -1168 289
rect -1202 187 -1168 221
rect -1202 119 -1168 153
rect -1202 51 -1168 85
rect -1202 -17 -1168 17
rect -1202 -85 -1168 -51
rect -1202 -153 -1168 -119
rect -1202 -221 -1168 -187
rect -1202 -289 -1168 -255
rect -1202 -357 -1168 -323
rect -1202 -425 -1168 -391
rect -1202 -493 -1168 -459
rect -1202 -561 -1168 -527
rect -1202 -629 -1168 -595
rect -1202 -697 -1168 -663
rect -1202 -765 -1168 -731
rect -1202 -833 -1168 -799
rect -1202 -901 -1168 -867
rect -1202 -969 -1168 -935
rect -1044 935 -1010 969
rect -1044 867 -1010 901
rect -1044 799 -1010 833
rect -1044 731 -1010 765
rect -1044 663 -1010 697
rect -1044 595 -1010 629
rect -1044 527 -1010 561
rect -1044 459 -1010 493
rect -1044 391 -1010 425
rect -1044 323 -1010 357
rect -1044 255 -1010 289
rect -1044 187 -1010 221
rect -1044 119 -1010 153
rect -1044 51 -1010 85
rect -1044 -17 -1010 17
rect -1044 -85 -1010 -51
rect -1044 -153 -1010 -119
rect -1044 -221 -1010 -187
rect -1044 -289 -1010 -255
rect -1044 -357 -1010 -323
rect -1044 -425 -1010 -391
rect -1044 -493 -1010 -459
rect -1044 -561 -1010 -527
rect -1044 -629 -1010 -595
rect -1044 -697 -1010 -663
rect -1044 -765 -1010 -731
rect -1044 -833 -1010 -799
rect -1044 -901 -1010 -867
rect -1044 -969 -1010 -935
rect -886 935 -852 969
rect -886 867 -852 901
rect -886 799 -852 833
rect -886 731 -852 765
rect -886 663 -852 697
rect -886 595 -852 629
rect -886 527 -852 561
rect -886 459 -852 493
rect -886 391 -852 425
rect -886 323 -852 357
rect -886 255 -852 289
rect -886 187 -852 221
rect -886 119 -852 153
rect -886 51 -852 85
rect -886 -17 -852 17
rect -886 -85 -852 -51
rect -886 -153 -852 -119
rect -886 -221 -852 -187
rect -886 -289 -852 -255
rect -886 -357 -852 -323
rect -886 -425 -852 -391
rect -886 -493 -852 -459
rect -886 -561 -852 -527
rect -886 -629 -852 -595
rect -886 -697 -852 -663
rect -886 -765 -852 -731
rect -886 -833 -852 -799
rect -886 -901 -852 -867
rect -886 -969 -852 -935
rect -728 935 -694 969
rect -728 867 -694 901
rect -728 799 -694 833
rect -728 731 -694 765
rect -728 663 -694 697
rect -728 595 -694 629
rect -728 527 -694 561
rect -728 459 -694 493
rect -728 391 -694 425
rect -728 323 -694 357
rect -728 255 -694 289
rect -728 187 -694 221
rect -728 119 -694 153
rect -728 51 -694 85
rect -728 -17 -694 17
rect -728 -85 -694 -51
rect -728 -153 -694 -119
rect -728 -221 -694 -187
rect -728 -289 -694 -255
rect -728 -357 -694 -323
rect -728 -425 -694 -391
rect -728 -493 -694 -459
rect -728 -561 -694 -527
rect -728 -629 -694 -595
rect -728 -697 -694 -663
rect -728 -765 -694 -731
rect -728 -833 -694 -799
rect -728 -901 -694 -867
rect -728 -969 -694 -935
rect -570 935 -536 969
rect -570 867 -536 901
rect -570 799 -536 833
rect -570 731 -536 765
rect -570 663 -536 697
rect -570 595 -536 629
rect -570 527 -536 561
rect -570 459 -536 493
rect -570 391 -536 425
rect -570 323 -536 357
rect -570 255 -536 289
rect -570 187 -536 221
rect -570 119 -536 153
rect -570 51 -536 85
rect -570 -17 -536 17
rect -570 -85 -536 -51
rect -570 -153 -536 -119
rect -570 -221 -536 -187
rect -570 -289 -536 -255
rect -570 -357 -536 -323
rect -570 -425 -536 -391
rect -570 -493 -536 -459
rect -570 -561 -536 -527
rect -570 -629 -536 -595
rect -570 -697 -536 -663
rect -570 -765 -536 -731
rect -570 -833 -536 -799
rect -570 -901 -536 -867
rect -570 -969 -536 -935
rect -412 935 -378 969
rect -412 867 -378 901
rect -412 799 -378 833
rect -412 731 -378 765
rect -412 663 -378 697
rect -412 595 -378 629
rect -412 527 -378 561
rect -412 459 -378 493
rect -412 391 -378 425
rect -412 323 -378 357
rect -412 255 -378 289
rect -412 187 -378 221
rect -412 119 -378 153
rect -412 51 -378 85
rect -412 -17 -378 17
rect -412 -85 -378 -51
rect -412 -153 -378 -119
rect -412 -221 -378 -187
rect -412 -289 -378 -255
rect -412 -357 -378 -323
rect -412 -425 -378 -391
rect -412 -493 -378 -459
rect -412 -561 -378 -527
rect -412 -629 -378 -595
rect -412 -697 -378 -663
rect -412 -765 -378 -731
rect -412 -833 -378 -799
rect -412 -901 -378 -867
rect -412 -969 -378 -935
rect -254 935 -220 969
rect -254 867 -220 901
rect -254 799 -220 833
rect -254 731 -220 765
rect -254 663 -220 697
rect -254 595 -220 629
rect -254 527 -220 561
rect -254 459 -220 493
rect -254 391 -220 425
rect -254 323 -220 357
rect -254 255 -220 289
rect -254 187 -220 221
rect -254 119 -220 153
rect -254 51 -220 85
rect -254 -17 -220 17
rect -254 -85 -220 -51
rect -254 -153 -220 -119
rect -254 -221 -220 -187
rect -254 -289 -220 -255
rect -254 -357 -220 -323
rect -254 -425 -220 -391
rect -254 -493 -220 -459
rect -254 -561 -220 -527
rect -254 -629 -220 -595
rect -254 -697 -220 -663
rect -254 -765 -220 -731
rect -254 -833 -220 -799
rect -254 -901 -220 -867
rect -254 -969 -220 -935
rect -96 935 -62 969
rect -96 867 -62 901
rect -96 799 -62 833
rect -96 731 -62 765
rect -96 663 -62 697
rect -96 595 -62 629
rect -96 527 -62 561
rect -96 459 -62 493
rect -96 391 -62 425
rect -96 323 -62 357
rect -96 255 -62 289
rect -96 187 -62 221
rect -96 119 -62 153
rect -96 51 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -51
rect -96 -153 -62 -119
rect -96 -221 -62 -187
rect -96 -289 -62 -255
rect -96 -357 -62 -323
rect -96 -425 -62 -391
rect -96 -493 -62 -459
rect -96 -561 -62 -527
rect -96 -629 -62 -595
rect -96 -697 -62 -663
rect -96 -765 -62 -731
rect -96 -833 -62 -799
rect -96 -901 -62 -867
rect -96 -969 -62 -935
rect 62 935 96 969
rect 62 867 96 901
rect 62 799 96 833
rect 62 731 96 765
rect 62 663 96 697
rect 62 595 96 629
rect 62 527 96 561
rect 62 459 96 493
rect 62 391 96 425
rect 62 323 96 357
rect 62 255 96 289
rect 62 187 96 221
rect 62 119 96 153
rect 62 51 96 85
rect 62 -17 96 17
rect 62 -85 96 -51
rect 62 -153 96 -119
rect 62 -221 96 -187
rect 62 -289 96 -255
rect 62 -357 96 -323
rect 62 -425 96 -391
rect 62 -493 96 -459
rect 62 -561 96 -527
rect 62 -629 96 -595
rect 62 -697 96 -663
rect 62 -765 96 -731
rect 62 -833 96 -799
rect 62 -901 96 -867
rect 62 -969 96 -935
rect 220 935 254 969
rect 220 867 254 901
rect 220 799 254 833
rect 220 731 254 765
rect 220 663 254 697
rect 220 595 254 629
rect 220 527 254 561
rect 220 459 254 493
rect 220 391 254 425
rect 220 323 254 357
rect 220 255 254 289
rect 220 187 254 221
rect 220 119 254 153
rect 220 51 254 85
rect 220 -17 254 17
rect 220 -85 254 -51
rect 220 -153 254 -119
rect 220 -221 254 -187
rect 220 -289 254 -255
rect 220 -357 254 -323
rect 220 -425 254 -391
rect 220 -493 254 -459
rect 220 -561 254 -527
rect 220 -629 254 -595
rect 220 -697 254 -663
rect 220 -765 254 -731
rect 220 -833 254 -799
rect 220 -901 254 -867
rect 220 -969 254 -935
rect 378 935 412 969
rect 378 867 412 901
rect 378 799 412 833
rect 378 731 412 765
rect 378 663 412 697
rect 378 595 412 629
rect 378 527 412 561
rect 378 459 412 493
rect 378 391 412 425
rect 378 323 412 357
rect 378 255 412 289
rect 378 187 412 221
rect 378 119 412 153
rect 378 51 412 85
rect 378 -17 412 17
rect 378 -85 412 -51
rect 378 -153 412 -119
rect 378 -221 412 -187
rect 378 -289 412 -255
rect 378 -357 412 -323
rect 378 -425 412 -391
rect 378 -493 412 -459
rect 378 -561 412 -527
rect 378 -629 412 -595
rect 378 -697 412 -663
rect 378 -765 412 -731
rect 378 -833 412 -799
rect 378 -901 412 -867
rect 378 -969 412 -935
rect 536 935 570 969
rect 536 867 570 901
rect 536 799 570 833
rect 536 731 570 765
rect 536 663 570 697
rect 536 595 570 629
rect 536 527 570 561
rect 536 459 570 493
rect 536 391 570 425
rect 536 323 570 357
rect 536 255 570 289
rect 536 187 570 221
rect 536 119 570 153
rect 536 51 570 85
rect 536 -17 570 17
rect 536 -85 570 -51
rect 536 -153 570 -119
rect 536 -221 570 -187
rect 536 -289 570 -255
rect 536 -357 570 -323
rect 536 -425 570 -391
rect 536 -493 570 -459
rect 536 -561 570 -527
rect 536 -629 570 -595
rect 536 -697 570 -663
rect 536 -765 570 -731
rect 536 -833 570 -799
rect 536 -901 570 -867
rect 536 -969 570 -935
rect 694 935 728 969
rect 694 867 728 901
rect 694 799 728 833
rect 694 731 728 765
rect 694 663 728 697
rect 694 595 728 629
rect 694 527 728 561
rect 694 459 728 493
rect 694 391 728 425
rect 694 323 728 357
rect 694 255 728 289
rect 694 187 728 221
rect 694 119 728 153
rect 694 51 728 85
rect 694 -17 728 17
rect 694 -85 728 -51
rect 694 -153 728 -119
rect 694 -221 728 -187
rect 694 -289 728 -255
rect 694 -357 728 -323
rect 694 -425 728 -391
rect 694 -493 728 -459
rect 694 -561 728 -527
rect 694 -629 728 -595
rect 694 -697 728 -663
rect 694 -765 728 -731
rect 694 -833 728 -799
rect 694 -901 728 -867
rect 694 -969 728 -935
rect 852 935 886 969
rect 852 867 886 901
rect 852 799 886 833
rect 852 731 886 765
rect 852 663 886 697
rect 852 595 886 629
rect 852 527 886 561
rect 852 459 886 493
rect 852 391 886 425
rect 852 323 886 357
rect 852 255 886 289
rect 852 187 886 221
rect 852 119 886 153
rect 852 51 886 85
rect 852 -17 886 17
rect 852 -85 886 -51
rect 852 -153 886 -119
rect 852 -221 886 -187
rect 852 -289 886 -255
rect 852 -357 886 -323
rect 852 -425 886 -391
rect 852 -493 886 -459
rect 852 -561 886 -527
rect 852 -629 886 -595
rect 852 -697 886 -663
rect 852 -765 886 -731
rect 852 -833 886 -799
rect 852 -901 886 -867
rect 852 -969 886 -935
rect 1010 935 1044 969
rect 1010 867 1044 901
rect 1010 799 1044 833
rect 1010 731 1044 765
rect 1010 663 1044 697
rect 1010 595 1044 629
rect 1010 527 1044 561
rect 1010 459 1044 493
rect 1010 391 1044 425
rect 1010 323 1044 357
rect 1010 255 1044 289
rect 1010 187 1044 221
rect 1010 119 1044 153
rect 1010 51 1044 85
rect 1010 -17 1044 17
rect 1010 -85 1044 -51
rect 1010 -153 1044 -119
rect 1010 -221 1044 -187
rect 1010 -289 1044 -255
rect 1010 -357 1044 -323
rect 1010 -425 1044 -391
rect 1010 -493 1044 -459
rect 1010 -561 1044 -527
rect 1010 -629 1044 -595
rect 1010 -697 1044 -663
rect 1010 -765 1044 -731
rect 1010 -833 1044 -799
rect 1010 -901 1044 -867
rect 1010 -969 1044 -935
rect 1168 935 1202 969
rect 1168 867 1202 901
rect 1168 799 1202 833
rect 1168 731 1202 765
rect 1168 663 1202 697
rect 1168 595 1202 629
rect 1168 527 1202 561
rect 1168 459 1202 493
rect 1168 391 1202 425
rect 1168 323 1202 357
rect 1168 255 1202 289
rect 1168 187 1202 221
rect 1168 119 1202 153
rect 1168 51 1202 85
rect 1168 -17 1202 17
rect 1168 -85 1202 -51
rect 1168 -153 1202 -119
rect 1168 -221 1202 -187
rect 1168 -289 1202 -255
rect 1168 -357 1202 -323
rect 1168 -425 1202 -391
rect 1168 -493 1202 -459
rect 1168 -561 1202 -527
rect 1168 -629 1202 -595
rect 1168 -697 1202 -663
rect 1168 -765 1202 -731
rect 1168 -833 1202 -799
rect 1168 -901 1202 -867
rect 1168 -969 1202 -935
<< nsubdiff >>
rect -1316 1149 -1207 1183
rect -1173 1149 -1139 1183
rect -1105 1149 -1071 1183
rect -1037 1149 -1003 1183
rect -969 1149 -935 1183
rect -901 1149 -867 1183
rect -833 1149 -799 1183
rect -765 1149 -731 1183
rect -697 1149 -663 1183
rect -629 1149 -595 1183
rect -561 1149 -527 1183
rect -493 1149 -459 1183
rect -425 1149 -391 1183
rect -357 1149 -323 1183
rect -289 1149 -255 1183
rect -221 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 221 1183
rect 255 1149 289 1183
rect 323 1149 357 1183
rect 391 1149 425 1183
rect 459 1149 493 1183
rect 527 1149 561 1183
rect 595 1149 629 1183
rect 663 1149 697 1183
rect 731 1149 765 1183
rect 799 1149 833 1183
rect 867 1149 901 1183
rect 935 1149 969 1183
rect 1003 1149 1037 1183
rect 1071 1149 1105 1183
rect 1139 1149 1173 1183
rect 1207 1149 1316 1183
rect -1316 1071 -1282 1149
rect -1316 1003 -1282 1037
rect 1282 1071 1316 1149
rect 1282 1003 1316 1037
rect -1316 935 -1282 969
rect -1316 867 -1282 901
rect -1316 799 -1282 833
rect -1316 731 -1282 765
rect -1316 663 -1282 697
rect -1316 595 -1282 629
rect -1316 527 -1282 561
rect -1316 459 -1282 493
rect -1316 391 -1282 425
rect -1316 323 -1282 357
rect -1316 255 -1282 289
rect -1316 187 -1282 221
rect -1316 119 -1282 153
rect -1316 51 -1282 85
rect -1316 -17 -1282 17
rect -1316 -85 -1282 -51
rect -1316 -153 -1282 -119
rect -1316 -221 -1282 -187
rect -1316 -289 -1282 -255
rect -1316 -357 -1282 -323
rect -1316 -425 -1282 -391
rect -1316 -493 -1282 -459
rect -1316 -561 -1282 -527
rect -1316 -629 -1282 -595
rect -1316 -697 -1282 -663
rect -1316 -765 -1282 -731
rect -1316 -833 -1282 -799
rect -1316 -901 -1282 -867
rect -1316 -969 -1282 -935
rect 1282 935 1316 969
rect 1282 867 1316 901
rect 1282 799 1316 833
rect 1282 731 1316 765
rect 1282 663 1316 697
rect 1282 595 1316 629
rect 1282 527 1316 561
rect 1282 459 1316 493
rect 1282 391 1316 425
rect 1282 323 1316 357
rect 1282 255 1316 289
rect 1282 187 1316 221
rect 1282 119 1316 153
rect 1282 51 1316 85
rect 1282 -17 1316 17
rect 1282 -85 1316 -51
rect 1282 -153 1316 -119
rect 1282 -221 1316 -187
rect 1282 -289 1316 -255
rect 1282 -357 1316 -323
rect 1282 -425 1316 -391
rect 1282 -493 1316 -459
rect 1282 -561 1316 -527
rect 1282 -629 1316 -595
rect 1282 -697 1316 -663
rect 1282 -765 1316 -731
rect 1282 -833 1316 -799
rect 1282 -901 1316 -867
rect 1282 -969 1316 -935
rect -1316 -1037 -1282 -1003
rect -1316 -1149 -1282 -1071
rect 1282 -1037 1316 -1003
rect 1282 -1149 1316 -1071
rect -1316 -1183 -1207 -1149
rect -1173 -1183 -1139 -1149
rect -1105 -1183 -1071 -1149
rect -1037 -1183 -1003 -1149
rect -969 -1183 -935 -1149
rect -901 -1183 -867 -1149
rect -833 -1183 -799 -1149
rect -765 -1183 -731 -1149
rect -697 -1183 -663 -1149
rect -629 -1183 -595 -1149
rect -561 -1183 -527 -1149
rect -493 -1183 -459 -1149
rect -425 -1183 -391 -1149
rect -357 -1183 -323 -1149
rect -289 -1183 -255 -1149
rect -221 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 221 -1149
rect 255 -1183 289 -1149
rect 323 -1183 357 -1149
rect 391 -1183 425 -1149
rect 459 -1183 493 -1149
rect 527 -1183 561 -1149
rect 595 -1183 629 -1149
rect 663 -1183 697 -1149
rect 731 -1183 765 -1149
rect 799 -1183 833 -1149
rect 867 -1183 901 -1149
rect 935 -1183 969 -1149
rect 1003 -1183 1037 -1149
rect 1071 -1183 1105 -1149
rect 1139 -1183 1173 -1149
rect 1207 -1183 1316 -1149
<< nsubdiffcont >>
rect -1207 1149 -1173 1183
rect -1139 1149 -1105 1183
rect -1071 1149 -1037 1183
rect -1003 1149 -969 1183
rect -935 1149 -901 1183
rect -867 1149 -833 1183
rect -799 1149 -765 1183
rect -731 1149 -697 1183
rect -663 1149 -629 1183
rect -595 1149 -561 1183
rect -527 1149 -493 1183
rect -459 1149 -425 1183
rect -391 1149 -357 1183
rect -323 1149 -289 1183
rect -255 1149 -221 1183
rect -187 1149 -153 1183
rect -119 1149 -85 1183
rect -51 1149 -17 1183
rect 17 1149 51 1183
rect 85 1149 119 1183
rect 153 1149 187 1183
rect 221 1149 255 1183
rect 289 1149 323 1183
rect 357 1149 391 1183
rect 425 1149 459 1183
rect 493 1149 527 1183
rect 561 1149 595 1183
rect 629 1149 663 1183
rect 697 1149 731 1183
rect 765 1149 799 1183
rect 833 1149 867 1183
rect 901 1149 935 1183
rect 969 1149 1003 1183
rect 1037 1149 1071 1183
rect 1105 1149 1139 1183
rect 1173 1149 1207 1183
rect -1316 1037 -1282 1071
rect -1316 969 -1282 1003
rect 1282 1037 1316 1071
rect -1316 901 -1282 935
rect -1316 833 -1282 867
rect -1316 765 -1282 799
rect -1316 697 -1282 731
rect -1316 629 -1282 663
rect -1316 561 -1282 595
rect -1316 493 -1282 527
rect -1316 425 -1282 459
rect -1316 357 -1282 391
rect -1316 289 -1282 323
rect -1316 221 -1282 255
rect -1316 153 -1282 187
rect -1316 85 -1282 119
rect -1316 17 -1282 51
rect -1316 -51 -1282 -17
rect -1316 -119 -1282 -85
rect -1316 -187 -1282 -153
rect -1316 -255 -1282 -221
rect -1316 -323 -1282 -289
rect -1316 -391 -1282 -357
rect -1316 -459 -1282 -425
rect -1316 -527 -1282 -493
rect -1316 -595 -1282 -561
rect -1316 -663 -1282 -629
rect -1316 -731 -1282 -697
rect -1316 -799 -1282 -765
rect -1316 -867 -1282 -833
rect -1316 -935 -1282 -901
rect -1316 -1003 -1282 -969
rect 1282 969 1316 1003
rect 1282 901 1316 935
rect 1282 833 1316 867
rect 1282 765 1316 799
rect 1282 697 1316 731
rect 1282 629 1316 663
rect 1282 561 1316 595
rect 1282 493 1316 527
rect 1282 425 1316 459
rect 1282 357 1316 391
rect 1282 289 1316 323
rect 1282 221 1316 255
rect 1282 153 1316 187
rect 1282 85 1316 119
rect 1282 17 1316 51
rect 1282 -51 1316 -17
rect 1282 -119 1316 -85
rect 1282 -187 1316 -153
rect 1282 -255 1316 -221
rect 1282 -323 1316 -289
rect 1282 -391 1316 -357
rect 1282 -459 1316 -425
rect 1282 -527 1316 -493
rect 1282 -595 1316 -561
rect 1282 -663 1316 -629
rect 1282 -731 1316 -697
rect 1282 -799 1316 -765
rect 1282 -867 1316 -833
rect 1282 -935 1316 -901
rect -1316 -1071 -1282 -1037
rect 1282 -1003 1316 -969
rect 1282 -1071 1316 -1037
rect -1207 -1183 -1173 -1149
rect -1139 -1183 -1105 -1149
rect -1071 -1183 -1037 -1149
rect -1003 -1183 -969 -1149
rect -935 -1183 -901 -1149
rect -867 -1183 -833 -1149
rect -799 -1183 -765 -1149
rect -731 -1183 -697 -1149
rect -663 -1183 -629 -1149
rect -595 -1183 -561 -1149
rect -527 -1183 -493 -1149
rect -459 -1183 -425 -1149
rect -391 -1183 -357 -1149
rect -323 -1183 -289 -1149
rect -255 -1183 -221 -1149
rect -187 -1183 -153 -1149
rect -119 -1183 -85 -1149
rect -51 -1183 -17 -1149
rect 17 -1183 51 -1149
rect 85 -1183 119 -1149
rect 153 -1183 187 -1149
rect 221 -1183 255 -1149
rect 289 -1183 323 -1149
rect 357 -1183 391 -1149
rect 425 -1183 459 -1149
rect 493 -1183 527 -1149
rect 561 -1183 595 -1149
rect 629 -1183 663 -1149
rect 697 -1183 731 -1149
rect 765 -1183 799 -1149
rect 833 -1183 867 -1149
rect 901 -1183 935 -1149
rect 969 -1183 1003 -1149
rect 1037 -1183 1071 -1149
rect 1105 -1183 1139 -1149
rect 1173 -1183 1207 -1149
<< poly >>
rect -1156 1081 -1056 1097
rect -1156 1047 -1123 1081
rect -1089 1047 -1056 1081
rect -1156 1000 -1056 1047
rect -998 1081 -898 1097
rect -998 1047 -965 1081
rect -931 1047 -898 1081
rect -998 1000 -898 1047
rect -840 1081 -740 1097
rect -840 1047 -807 1081
rect -773 1047 -740 1081
rect -840 1000 -740 1047
rect -682 1081 -582 1097
rect -682 1047 -649 1081
rect -615 1047 -582 1081
rect -682 1000 -582 1047
rect -524 1081 -424 1097
rect -524 1047 -491 1081
rect -457 1047 -424 1081
rect -524 1000 -424 1047
rect -366 1081 -266 1097
rect -366 1047 -333 1081
rect -299 1047 -266 1081
rect -366 1000 -266 1047
rect -208 1081 -108 1097
rect -208 1047 -175 1081
rect -141 1047 -108 1081
rect -208 1000 -108 1047
rect -50 1081 50 1097
rect -50 1047 -17 1081
rect 17 1047 50 1081
rect -50 1000 50 1047
rect 108 1081 208 1097
rect 108 1047 141 1081
rect 175 1047 208 1081
rect 108 1000 208 1047
rect 266 1081 366 1097
rect 266 1047 299 1081
rect 333 1047 366 1081
rect 266 1000 366 1047
rect 424 1081 524 1097
rect 424 1047 457 1081
rect 491 1047 524 1081
rect 424 1000 524 1047
rect 582 1081 682 1097
rect 582 1047 615 1081
rect 649 1047 682 1081
rect 582 1000 682 1047
rect 740 1081 840 1097
rect 740 1047 773 1081
rect 807 1047 840 1081
rect 740 1000 840 1047
rect 898 1081 998 1097
rect 898 1047 931 1081
rect 965 1047 998 1081
rect 898 1000 998 1047
rect 1056 1081 1156 1097
rect 1056 1047 1089 1081
rect 1123 1047 1156 1081
rect 1056 1000 1156 1047
rect -1156 -1047 -1056 -1000
rect -1156 -1081 -1123 -1047
rect -1089 -1081 -1056 -1047
rect -1156 -1097 -1056 -1081
rect -998 -1047 -898 -1000
rect -998 -1081 -965 -1047
rect -931 -1081 -898 -1047
rect -998 -1097 -898 -1081
rect -840 -1047 -740 -1000
rect -840 -1081 -807 -1047
rect -773 -1081 -740 -1047
rect -840 -1097 -740 -1081
rect -682 -1047 -582 -1000
rect -682 -1081 -649 -1047
rect -615 -1081 -582 -1047
rect -682 -1097 -582 -1081
rect -524 -1047 -424 -1000
rect -524 -1081 -491 -1047
rect -457 -1081 -424 -1047
rect -524 -1097 -424 -1081
rect -366 -1047 -266 -1000
rect -366 -1081 -333 -1047
rect -299 -1081 -266 -1047
rect -366 -1097 -266 -1081
rect -208 -1047 -108 -1000
rect -208 -1081 -175 -1047
rect -141 -1081 -108 -1047
rect -208 -1097 -108 -1081
rect -50 -1047 50 -1000
rect -50 -1081 -17 -1047
rect 17 -1081 50 -1047
rect -50 -1097 50 -1081
rect 108 -1047 208 -1000
rect 108 -1081 141 -1047
rect 175 -1081 208 -1047
rect 108 -1097 208 -1081
rect 266 -1047 366 -1000
rect 266 -1081 299 -1047
rect 333 -1081 366 -1047
rect 266 -1097 366 -1081
rect 424 -1047 524 -1000
rect 424 -1081 457 -1047
rect 491 -1081 524 -1047
rect 424 -1097 524 -1081
rect 582 -1047 682 -1000
rect 582 -1081 615 -1047
rect 649 -1081 682 -1047
rect 582 -1097 682 -1081
rect 740 -1047 840 -1000
rect 740 -1081 773 -1047
rect 807 -1081 840 -1047
rect 740 -1097 840 -1081
rect 898 -1047 998 -1000
rect 898 -1081 931 -1047
rect 965 -1081 998 -1047
rect 898 -1097 998 -1081
rect 1056 -1047 1156 -1000
rect 1056 -1081 1089 -1047
rect 1123 -1081 1156 -1047
rect 1056 -1097 1156 -1081
<< polycont >>
rect -1123 1047 -1089 1081
rect -965 1047 -931 1081
rect -807 1047 -773 1081
rect -649 1047 -615 1081
rect -491 1047 -457 1081
rect -333 1047 -299 1081
rect -175 1047 -141 1081
rect -17 1047 17 1081
rect 141 1047 175 1081
rect 299 1047 333 1081
rect 457 1047 491 1081
rect 615 1047 649 1081
rect 773 1047 807 1081
rect 931 1047 965 1081
rect 1089 1047 1123 1081
rect -1123 -1081 -1089 -1047
rect -965 -1081 -931 -1047
rect -807 -1081 -773 -1047
rect -649 -1081 -615 -1047
rect -491 -1081 -457 -1047
rect -333 -1081 -299 -1047
rect -175 -1081 -141 -1047
rect -17 -1081 17 -1047
rect 141 -1081 175 -1047
rect 299 -1081 333 -1047
rect 457 -1081 491 -1047
rect 615 -1081 649 -1047
rect 773 -1081 807 -1047
rect 931 -1081 965 -1047
rect 1089 -1081 1123 -1047
<< locali >>
rect -1316 1149 -1207 1183
rect -1173 1149 -1139 1183
rect -1105 1149 -1071 1183
rect -1037 1149 -1003 1183
rect -969 1149 -935 1183
rect -901 1149 -867 1183
rect -833 1149 -799 1183
rect -765 1149 -731 1183
rect -697 1149 -663 1183
rect -629 1149 -595 1183
rect -561 1149 -527 1183
rect -493 1149 -459 1183
rect -425 1149 -391 1183
rect -357 1149 -323 1183
rect -289 1149 -255 1183
rect -221 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 221 1183
rect 255 1149 289 1183
rect 323 1149 357 1183
rect 391 1149 425 1183
rect 459 1149 493 1183
rect 527 1149 561 1183
rect 595 1149 629 1183
rect 663 1149 697 1183
rect 731 1149 765 1183
rect 799 1149 833 1183
rect 867 1149 901 1183
rect 935 1149 969 1183
rect 1003 1149 1037 1183
rect 1071 1149 1105 1183
rect 1139 1149 1173 1183
rect 1207 1149 1316 1183
rect -1316 1071 -1282 1149
rect -1156 1047 -1123 1081
rect -1089 1047 -1056 1081
rect -998 1047 -965 1081
rect -931 1047 -898 1081
rect -840 1047 -807 1081
rect -773 1047 -740 1081
rect -682 1047 -649 1081
rect -615 1047 -582 1081
rect -524 1047 -491 1081
rect -457 1047 -424 1081
rect -366 1047 -333 1081
rect -299 1047 -266 1081
rect -208 1047 -175 1081
rect -141 1047 -108 1081
rect -50 1047 -17 1081
rect 17 1047 50 1081
rect 108 1047 141 1081
rect 175 1047 208 1081
rect 266 1047 299 1081
rect 333 1047 366 1081
rect 424 1047 457 1081
rect 491 1047 524 1081
rect 582 1047 615 1081
rect 649 1047 682 1081
rect 740 1047 773 1081
rect 807 1047 840 1081
rect 898 1047 931 1081
rect 965 1047 998 1081
rect 1056 1047 1089 1081
rect 1123 1047 1156 1081
rect 1282 1071 1316 1149
rect -1316 1003 -1282 1037
rect -1316 935 -1282 969
rect -1316 867 -1282 901
rect -1316 799 -1282 833
rect -1316 731 -1282 765
rect -1316 663 -1282 697
rect -1316 595 -1282 629
rect -1316 527 -1282 561
rect -1316 459 -1282 493
rect -1316 391 -1282 425
rect -1316 323 -1282 357
rect -1316 255 -1282 289
rect -1316 187 -1282 221
rect -1316 119 -1282 153
rect -1316 51 -1282 85
rect -1316 -17 -1282 17
rect -1316 -85 -1282 -51
rect -1316 -153 -1282 -119
rect -1316 -221 -1282 -187
rect -1316 -289 -1282 -255
rect -1316 -357 -1282 -323
rect -1316 -425 -1282 -391
rect -1316 -493 -1282 -459
rect -1316 -561 -1282 -527
rect -1316 -629 -1282 -595
rect -1316 -697 -1282 -663
rect -1316 -765 -1282 -731
rect -1316 -833 -1282 -799
rect -1316 -901 -1282 -867
rect -1316 -969 -1282 -935
rect -1316 -1037 -1282 -1003
rect -1202 969 -1168 1004
rect -1202 901 -1168 935
rect -1202 833 -1168 867
rect -1202 765 -1168 799
rect -1202 697 -1168 731
rect -1202 629 -1168 663
rect -1202 561 -1168 595
rect -1202 493 -1168 527
rect -1202 425 -1168 459
rect -1202 357 -1168 391
rect -1202 289 -1168 323
rect -1202 221 -1168 255
rect -1202 153 -1168 187
rect -1202 85 -1168 119
rect -1202 17 -1168 51
rect -1202 -51 -1168 -17
rect -1202 -119 -1168 -85
rect -1202 -187 -1168 -153
rect -1202 -255 -1168 -221
rect -1202 -323 -1168 -289
rect -1202 -391 -1168 -357
rect -1202 -459 -1168 -425
rect -1202 -527 -1168 -493
rect -1202 -595 -1168 -561
rect -1202 -663 -1168 -629
rect -1202 -731 -1168 -697
rect -1202 -799 -1168 -765
rect -1202 -867 -1168 -833
rect -1202 -935 -1168 -901
rect -1202 -1004 -1168 -969
rect -1044 969 -1010 1004
rect -1044 901 -1010 935
rect -1044 833 -1010 867
rect -1044 765 -1010 799
rect -1044 697 -1010 731
rect -1044 629 -1010 663
rect -1044 561 -1010 595
rect -1044 493 -1010 527
rect -1044 425 -1010 459
rect -1044 357 -1010 391
rect -1044 289 -1010 323
rect -1044 221 -1010 255
rect -1044 153 -1010 187
rect -1044 85 -1010 119
rect -1044 17 -1010 51
rect -1044 -51 -1010 -17
rect -1044 -119 -1010 -85
rect -1044 -187 -1010 -153
rect -1044 -255 -1010 -221
rect -1044 -323 -1010 -289
rect -1044 -391 -1010 -357
rect -1044 -459 -1010 -425
rect -1044 -527 -1010 -493
rect -1044 -595 -1010 -561
rect -1044 -663 -1010 -629
rect -1044 -731 -1010 -697
rect -1044 -799 -1010 -765
rect -1044 -867 -1010 -833
rect -1044 -935 -1010 -901
rect -1044 -1004 -1010 -969
rect -886 969 -852 1004
rect -886 901 -852 935
rect -886 833 -852 867
rect -886 765 -852 799
rect -886 697 -852 731
rect -886 629 -852 663
rect -886 561 -852 595
rect -886 493 -852 527
rect -886 425 -852 459
rect -886 357 -852 391
rect -886 289 -852 323
rect -886 221 -852 255
rect -886 153 -852 187
rect -886 85 -852 119
rect -886 17 -852 51
rect -886 -51 -852 -17
rect -886 -119 -852 -85
rect -886 -187 -852 -153
rect -886 -255 -852 -221
rect -886 -323 -852 -289
rect -886 -391 -852 -357
rect -886 -459 -852 -425
rect -886 -527 -852 -493
rect -886 -595 -852 -561
rect -886 -663 -852 -629
rect -886 -731 -852 -697
rect -886 -799 -852 -765
rect -886 -867 -852 -833
rect -886 -935 -852 -901
rect -886 -1004 -852 -969
rect -728 969 -694 1004
rect -728 901 -694 935
rect -728 833 -694 867
rect -728 765 -694 799
rect -728 697 -694 731
rect -728 629 -694 663
rect -728 561 -694 595
rect -728 493 -694 527
rect -728 425 -694 459
rect -728 357 -694 391
rect -728 289 -694 323
rect -728 221 -694 255
rect -728 153 -694 187
rect -728 85 -694 119
rect -728 17 -694 51
rect -728 -51 -694 -17
rect -728 -119 -694 -85
rect -728 -187 -694 -153
rect -728 -255 -694 -221
rect -728 -323 -694 -289
rect -728 -391 -694 -357
rect -728 -459 -694 -425
rect -728 -527 -694 -493
rect -728 -595 -694 -561
rect -728 -663 -694 -629
rect -728 -731 -694 -697
rect -728 -799 -694 -765
rect -728 -867 -694 -833
rect -728 -935 -694 -901
rect -728 -1004 -694 -969
rect -570 969 -536 1004
rect -570 901 -536 935
rect -570 833 -536 867
rect -570 765 -536 799
rect -570 697 -536 731
rect -570 629 -536 663
rect -570 561 -536 595
rect -570 493 -536 527
rect -570 425 -536 459
rect -570 357 -536 391
rect -570 289 -536 323
rect -570 221 -536 255
rect -570 153 -536 187
rect -570 85 -536 119
rect -570 17 -536 51
rect -570 -51 -536 -17
rect -570 -119 -536 -85
rect -570 -187 -536 -153
rect -570 -255 -536 -221
rect -570 -323 -536 -289
rect -570 -391 -536 -357
rect -570 -459 -536 -425
rect -570 -527 -536 -493
rect -570 -595 -536 -561
rect -570 -663 -536 -629
rect -570 -731 -536 -697
rect -570 -799 -536 -765
rect -570 -867 -536 -833
rect -570 -935 -536 -901
rect -570 -1004 -536 -969
rect -412 969 -378 1004
rect -412 901 -378 935
rect -412 833 -378 867
rect -412 765 -378 799
rect -412 697 -378 731
rect -412 629 -378 663
rect -412 561 -378 595
rect -412 493 -378 527
rect -412 425 -378 459
rect -412 357 -378 391
rect -412 289 -378 323
rect -412 221 -378 255
rect -412 153 -378 187
rect -412 85 -378 119
rect -412 17 -378 51
rect -412 -51 -378 -17
rect -412 -119 -378 -85
rect -412 -187 -378 -153
rect -412 -255 -378 -221
rect -412 -323 -378 -289
rect -412 -391 -378 -357
rect -412 -459 -378 -425
rect -412 -527 -378 -493
rect -412 -595 -378 -561
rect -412 -663 -378 -629
rect -412 -731 -378 -697
rect -412 -799 -378 -765
rect -412 -867 -378 -833
rect -412 -935 -378 -901
rect -412 -1004 -378 -969
rect -254 969 -220 1004
rect -254 901 -220 935
rect -254 833 -220 867
rect -254 765 -220 799
rect -254 697 -220 731
rect -254 629 -220 663
rect -254 561 -220 595
rect -254 493 -220 527
rect -254 425 -220 459
rect -254 357 -220 391
rect -254 289 -220 323
rect -254 221 -220 255
rect -254 153 -220 187
rect -254 85 -220 119
rect -254 17 -220 51
rect -254 -51 -220 -17
rect -254 -119 -220 -85
rect -254 -187 -220 -153
rect -254 -255 -220 -221
rect -254 -323 -220 -289
rect -254 -391 -220 -357
rect -254 -459 -220 -425
rect -254 -527 -220 -493
rect -254 -595 -220 -561
rect -254 -663 -220 -629
rect -254 -731 -220 -697
rect -254 -799 -220 -765
rect -254 -867 -220 -833
rect -254 -935 -220 -901
rect -254 -1004 -220 -969
rect -96 969 -62 1004
rect -96 901 -62 935
rect -96 833 -62 867
rect -96 765 -62 799
rect -96 697 -62 731
rect -96 629 -62 663
rect -96 561 -62 595
rect -96 493 -62 527
rect -96 425 -62 459
rect -96 357 -62 391
rect -96 289 -62 323
rect -96 221 -62 255
rect -96 153 -62 187
rect -96 85 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -85
rect -96 -187 -62 -153
rect -96 -255 -62 -221
rect -96 -323 -62 -289
rect -96 -391 -62 -357
rect -96 -459 -62 -425
rect -96 -527 -62 -493
rect -96 -595 -62 -561
rect -96 -663 -62 -629
rect -96 -731 -62 -697
rect -96 -799 -62 -765
rect -96 -867 -62 -833
rect -96 -935 -62 -901
rect -96 -1004 -62 -969
rect 62 969 96 1004
rect 62 901 96 935
rect 62 833 96 867
rect 62 765 96 799
rect 62 697 96 731
rect 62 629 96 663
rect 62 561 96 595
rect 62 493 96 527
rect 62 425 96 459
rect 62 357 96 391
rect 62 289 96 323
rect 62 221 96 255
rect 62 153 96 187
rect 62 85 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -85
rect 62 -187 96 -153
rect 62 -255 96 -221
rect 62 -323 96 -289
rect 62 -391 96 -357
rect 62 -459 96 -425
rect 62 -527 96 -493
rect 62 -595 96 -561
rect 62 -663 96 -629
rect 62 -731 96 -697
rect 62 -799 96 -765
rect 62 -867 96 -833
rect 62 -935 96 -901
rect 62 -1004 96 -969
rect 220 969 254 1004
rect 220 901 254 935
rect 220 833 254 867
rect 220 765 254 799
rect 220 697 254 731
rect 220 629 254 663
rect 220 561 254 595
rect 220 493 254 527
rect 220 425 254 459
rect 220 357 254 391
rect 220 289 254 323
rect 220 221 254 255
rect 220 153 254 187
rect 220 85 254 119
rect 220 17 254 51
rect 220 -51 254 -17
rect 220 -119 254 -85
rect 220 -187 254 -153
rect 220 -255 254 -221
rect 220 -323 254 -289
rect 220 -391 254 -357
rect 220 -459 254 -425
rect 220 -527 254 -493
rect 220 -595 254 -561
rect 220 -663 254 -629
rect 220 -731 254 -697
rect 220 -799 254 -765
rect 220 -867 254 -833
rect 220 -935 254 -901
rect 220 -1004 254 -969
rect 378 969 412 1004
rect 378 901 412 935
rect 378 833 412 867
rect 378 765 412 799
rect 378 697 412 731
rect 378 629 412 663
rect 378 561 412 595
rect 378 493 412 527
rect 378 425 412 459
rect 378 357 412 391
rect 378 289 412 323
rect 378 221 412 255
rect 378 153 412 187
rect 378 85 412 119
rect 378 17 412 51
rect 378 -51 412 -17
rect 378 -119 412 -85
rect 378 -187 412 -153
rect 378 -255 412 -221
rect 378 -323 412 -289
rect 378 -391 412 -357
rect 378 -459 412 -425
rect 378 -527 412 -493
rect 378 -595 412 -561
rect 378 -663 412 -629
rect 378 -731 412 -697
rect 378 -799 412 -765
rect 378 -867 412 -833
rect 378 -935 412 -901
rect 378 -1004 412 -969
rect 536 969 570 1004
rect 536 901 570 935
rect 536 833 570 867
rect 536 765 570 799
rect 536 697 570 731
rect 536 629 570 663
rect 536 561 570 595
rect 536 493 570 527
rect 536 425 570 459
rect 536 357 570 391
rect 536 289 570 323
rect 536 221 570 255
rect 536 153 570 187
rect 536 85 570 119
rect 536 17 570 51
rect 536 -51 570 -17
rect 536 -119 570 -85
rect 536 -187 570 -153
rect 536 -255 570 -221
rect 536 -323 570 -289
rect 536 -391 570 -357
rect 536 -459 570 -425
rect 536 -527 570 -493
rect 536 -595 570 -561
rect 536 -663 570 -629
rect 536 -731 570 -697
rect 536 -799 570 -765
rect 536 -867 570 -833
rect 536 -935 570 -901
rect 536 -1004 570 -969
rect 694 969 728 1004
rect 694 901 728 935
rect 694 833 728 867
rect 694 765 728 799
rect 694 697 728 731
rect 694 629 728 663
rect 694 561 728 595
rect 694 493 728 527
rect 694 425 728 459
rect 694 357 728 391
rect 694 289 728 323
rect 694 221 728 255
rect 694 153 728 187
rect 694 85 728 119
rect 694 17 728 51
rect 694 -51 728 -17
rect 694 -119 728 -85
rect 694 -187 728 -153
rect 694 -255 728 -221
rect 694 -323 728 -289
rect 694 -391 728 -357
rect 694 -459 728 -425
rect 694 -527 728 -493
rect 694 -595 728 -561
rect 694 -663 728 -629
rect 694 -731 728 -697
rect 694 -799 728 -765
rect 694 -867 728 -833
rect 694 -935 728 -901
rect 694 -1004 728 -969
rect 852 969 886 1004
rect 852 901 886 935
rect 852 833 886 867
rect 852 765 886 799
rect 852 697 886 731
rect 852 629 886 663
rect 852 561 886 595
rect 852 493 886 527
rect 852 425 886 459
rect 852 357 886 391
rect 852 289 886 323
rect 852 221 886 255
rect 852 153 886 187
rect 852 85 886 119
rect 852 17 886 51
rect 852 -51 886 -17
rect 852 -119 886 -85
rect 852 -187 886 -153
rect 852 -255 886 -221
rect 852 -323 886 -289
rect 852 -391 886 -357
rect 852 -459 886 -425
rect 852 -527 886 -493
rect 852 -595 886 -561
rect 852 -663 886 -629
rect 852 -731 886 -697
rect 852 -799 886 -765
rect 852 -867 886 -833
rect 852 -935 886 -901
rect 852 -1004 886 -969
rect 1010 969 1044 1004
rect 1010 901 1044 935
rect 1010 833 1044 867
rect 1010 765 1044 799
rect 1010 697 1044 731
rect 1010 629 1044 663
rect 1010 561 1044 595
rect 1010 493 1044 527
rect 1010 425 1044 459
rect 1010 357 1044 391
rect 1010 289 1044 323
rect 1010 221 1044 255
rect 1010 153 1044 187
rect 1010 85 1044 119
rect 1010 17 1044 51
rect 1010 -51 1044 -17
rect 1010 -119 1044 -85
rect 1010 -187 1044 -153
rect 1010 -255 1044 -221
rect 1010 -323 1044 -289
rect 1010 -391 1044 -357
rect 1010 -459 1044 -425
rect 1010 -527 1044 -493
rect 1010 -595 1044 -561
rect 1010 -663 1044 -629
rect 1010 -731 1044 -697
rect 1010 -799 1044 -765
rect 1010 -867 1044 -833
rect 1010 -935 1044 -901
rect 1010 -1004 1044 -969
rect 1168 969 1202 1004
rect 1168 901 1202 935
rect 1168 833 1202 867
rect 1168 765 1202 799
rect 1168 697 1202 731
rect 1168 629 1202 663
rect 1168 561 1202 595
rect 1168 493 1202 527
rect 1168 425 1202 459
rect 1168 357 1202 391
rect 1168 289 1202 323
rect 1168 221 1202 255
rect 1168 153 1202 187
rect 1168 85 1202 119
rect 1168 17 1202 51
rect 1168 -51 1202 -17
rect 1168 -119 1202 -85
rect 1168 -187 1202 -153
rect 1168 -255 1202 -221
rect 1168 -323 1202 -289
rect 1168 -391 1202 -357
rect 1168 -459 1202 -425
rect 1168 -527 1202 -493
rect 1168 -595 1202 -561
rect 1168 -663 1202 -629
rect 1168 -731 1202 -697
rect 1168 -799 1202 -765
rect 1168 -867 1202 -833
rect 1168 -935 1202 -901
rect 1168 -1004 1202 -969
rect 1282 1003 1316 1037
rect 1282 935 1316 969
rect 1282 867 1316 901
rect 1282 799 1316 833
rect 1282 731 1316 765
rect 1282 663 1316 697
rect 1282 595 1316 629
rect 1282 527 1316 561
rect 1282 459 1316 493
rect 1282 391 1316 425
rect 1282 323 1316 357
rect 1282 255 1316 289
rect 1282 187 1316 221
rect 1282 119 1316 153
rect 1282 51 1316 85
rect 1282 -17 1316 17
rect 1282 -85 1316 -51
rect 1282 -153 1316 -119
rect 1282 -221 1316 -187
rect 1282 -289 1316 -255
rect 1282 -357 1316 -323
rect 1282 -425 1316 -391
rect 1282 -493 1316 -459
rect 1282 -561 1316 -527
rect 1282 -629 1316 -595
rect 1282 -697 1316 -663
rect 1282 -765 1316 -731
rect 1282 -833 1316 -799
rect 1282 -901 1316 -867
rect 1282 -969 1316 -935
rect 1282 -1037 1316 -1003
rect -1316 -1149 -1282 -1071
rect -1156 -1081 -1123 -1047
rect -1089 -1081 -1056 -1047
rect -998 -1081 -965 -1047
rect -931 -1081 -898 -1047
rect -840 -1081 -807 -1047
rect -773 -1081 -740 -1047
rect -682 -1081 -649 -1047
rect -615 -1081 -582 -1047
rect -524 -1081 -491 -1047
rect -457 -1081 -424 -1047
rect -366 -1081 -333 -1047
rect -299 -1081 -266 -1047
rect -208 -1081 -175 -1047
rect -141 -1081 -108 -1047
rect -50 -1081 -17 -1047
rect 17 -1081 50 -1047
rect 108 -1081 141 -1047
rect 175 -1081 208 -1047
rect 266 -1081 299 -1047
rect 333 -1081 366 -1047
rect 424 -1081 457 -1047
rect 491 -1081 524 -1047
rect 582 -1081 615 -1047
rect 649 -1081 682 -1047
rect 740 -1081 773 -1047
rect 807 -1081 840 -1047
rect 898 -1081 931 -1047
rect 965 -1081 998 -1047
rect 1056 -1081 1089 -1047
rect 1123 -1081 1156 -1047
rect 1282 -1149 1316 -1071
rect -1316 -1183 -1207 -1149
rect -1173 -1183 -1139 -1149
rect -1105 -1183 -1071 -1149
rect -1037 -1183 -1003 -1149
rect -969 -1183 -935 -1149
rect -901 -1183 -867 -1149
rect -833 -1183 -799 -1149
rect -765 -1183 -731 -1149
rect -697 -1183 -663 -1149
rect -629 -1183 -595 -1149
rect -561 -1183 -527 -1149
rect -493 -1183 -459 -1149
rect -425 -1183 -391 -1149
rect -357 -1183 -323 -1149
rect -289 -1183 -255 -1149
rect -221 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 221 -1149
rect 255 -1183 289 -1149
rect 323 -1183 357 -1149
rect 391 -1183 425 -1149
rect 459 -1183 493 -1149
rect 527 -1183 561 -1149
rect 595 -1183 629 -1149
rect 663 -1183 697 -1149
rect 731 -1183 765 -1149
rect 799 -1183 833 -1149
rect 867 -1183 901 -1149
rect 935 -1183 969 -1149
rect 1003 -1183 1037 -1149
rect 1071 -1183 1105 -1149
rect 1139 -1183 1173 -1149
rect 1207 -1183 1316 -1149
<< properties >>
string FIXED_BBOX -1299 -1166 1299 1166
<< end >>
