magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< pwell >>
rect -324 1628 324 1662
rect -324 -1628 -290 1628
rect 290 -1628 324 1628
rect -324 -1662 324 -1628
<< psubdiff >>
rect -324 1628 -221 1662
rect -187 1628 -153 1662
rect -119 1628 -85 1662
rect -51 1628 -17 1662
rect 17 1628 51 1662
rect 85 1628 119 1662
rect 153 1628 187 1662
rect 221 1628 324 1662
rect -324 1547 -290 1628
rect 290 1547 324 1628
rect -324 1479 -290 1513
rect -324 1411 -290 1445
rect -324 1343 -290 1377
rect -324 1275 -290 1309
rect -324 1207 -290 1241
rect -324 1139 -290 1173
rect -324 1071 -290 1105
rect -324 1003 -290 1037
rect -324 935 -290 969
rect -324 867 -290 901
rect -324 799 -290 833
rect -324 731 -290 765
rect -324 663 -290 697
rect -324 595 -290 629
rect -324 527 -290 561
rect -324 459 -290 493
rect -324 391 -290 425
rect -324 323 -290 357
rect -324 255 -290 289
rect -324 187 -290 221
rect -324 119 -290 153
rect -324 51 -290 85
rect -324 -17 -290 17
rect -324 -85 -290 -51
rect -324 -153 -290 -119
rect -324 -221 -290 -187
rect -324 -289 -290 -255
rect -324 -357 -290 -323
rect -324 -425 -290 -391
rect -324 -493 -290 -459
rect -324 -561 -290 -527
rect -324 -629 -290 -595
rect -324 -697 -290 -663
rect -324 -765 -290 -731
rect -324 -833 -290 -799
rect -324 -901 -290 -867
rect -324 -969 -290 -935
rect -324 -1037 -290 -1003
rect -324 -1105 -290 -1071
rect -324 -1173 -290 -1139
rect -324 -1241 -290 -1207
rect -324 -1309 -290 -1275
rect -324 -1377 -290 -1343
rect -324 -1445 -290 -1411
rect -324 -1513 -290 -1479
rect 290 1479 324 1513
rect 290 1411 324 1445
rect 290 1343 324 1377
rect 290 1275 324 1309
rect 290 1207 324 1241
rect 290 1139 324 1173
rect 290 1071 324 1105
rect 290 1003 324 1037
rect 290 935 324 969
rect 290 867 324 901
rect 290 799 324 833
rect 290 731 324 765
rect 290 663 324 697
rect 290 595 324 629
rect 290 527 324 561
rect 290 459 324 493
rect 290 391 324 425
rect 290 323 324 357
rect 290 255 324 289
rect 290 187 324 221
rect 290 119 324 153
rect 290 51 324 85
rect 290 -17 324 17
rect 290 -85 324 -51
rect 290 -153 324 -119
rect 290 -221 324 -187
rect 290 -289 324 -255
rect 290 -357 324 -323
rect 290 -425 324 -391
rect 290 -493 324 -459
rect 290 -561 324 -527
rect 290 -629 324 -595
rect 290 -697 324 -663
rect 290 -765 324 -731
rect 290 -833 324 -799
rect 290 -901 324 -867
rect 290 -969 324 -935
rect 290 -1037 324 -1003
rect 290 -1105 324 -1071
rect 290 -1173 324 -1139
rect 290 -1241 324 -1207
rect 290 -1309 324 -1275
rect 290 -1377 324 -1343
rect 290 -1445 324 -1411
rect 290 -1513 324 -1479
rect -324 -1628 -290 -1547
rect 290 -1628 324 -1547
rect -324 -1662 -221 -1628
rect -187 -1662 -153 -1628
rect -119 -1662 -85 -1628
rect -51 -1662 -17 -1628
rect 17 -1662 51 -1628
rect 85 -1662 119 -1628
rect 153 -1662 187 -1628
rect 221 -1662 324 -1628
<< psubdiffcont >>
rect -221 1628 -187 1662
rect -153 1628 -119 1662
rect -85 1628 -51 1662
rect -17 1628 17 1662
rect 51 1628 85 1662
rect 119 1628 153 1662
rect 187 1628 221 1662
rect -324 1513 -290 1547
rect -324 1445 -290 1479
rect -324 1377 -290 1411
rect -324 1309 -290 1343
rect -324 1241 -290 1275
rect -324 1173 -290 1207
rect -324 1105 -290 1139
rect -324 1037 -290 1071
rect -324 969 -290 1003
rect -324 901 -290 935
rect -324 833 -290 867
rect -324 765 -290 799
rect -324 697 -290 731
rect -324 629 -290 663
rect -324 561 -290 595
rect -324 493 -290 527
rect -324 425 -290 459
rect -324 357 -290 391
rect -324 289 -290 323
rect -324 221 -290 255
rect -324 153 -290 187
rect -324 85 -290 119
rect -324 17 -290 51
rect -324 -51 -290 -17
rect -324 -119 -290 -85
rect -324 -187 -290 -153
rect -324 -255 -290 -221
rect -324 -323 -290 -289
rect -324 -391 -290 -357
rect -324 -459 -290 -425
rect -324 -527 -290 -493
rect -324 -595 -290 -561
rect -324 -663 -290 -629
rect -324 -731 -290 -697
rect -324 -799 -290 -765
rect -324 -867 -290 -833
rect -324 -935 -290 -901
rect -324 -1003 -290 -969
rect -324 -1071 -290 -1037
rect -324 -1139 -290 -1105
rect -324 -1207 -290 -1173
rect -324 -1275 -290 -1241
rect -324 -1343 -290 -1309
rect -324 -1411 -290 -1377
rect -324 -1479 -290 -1445
rect -324 -1547 -290 -1513
rect 290 1513 324 1547
rect 290 1445 324 1479
rect 290 1377 324 1411
rect 290 1309 324 1343
rect 290 1241 324 1275
rect 290 1173 324 1207
rect 290 1105 324 1139
rect 290 1037 324 1071
rect 290 969 324 1003
rect 290 901 324 935
rect 290 833 324 867
rect 290 765 324 799
rect 290 697 324 731
rect 290 629 324 663
rect 290 561 324 595
rect 290 493 324 527
rect 290 425 324 459
rect 290 357 324 391
rect 290 289 324 323
rect 290 221 324 255
rect 290 153 324 187
rect 290 85 324 119
rect 290 17 324 51
rect 290 -51 324 -17
rect 290 -119 324 -85
rect 290 -187 324 -153
rect 290 -255 324 -221
rect 290 -323 324 -289
rect 290 -391 324 -357
rect 290 -459 324 -425
rect 290 -527 324 -493
rect 290 -595 324 -561
rect 290 -663 324 -629
rect 290 -731 324 -697
rect 290 -799 324 -765
rect 290 -867 324 -833
rect 290 -935 324 -901
rect 290 -1003 324 -969
rect 290 -1071 324 -1037
rect 290 -1139 324 -1105
rect 290 -1207 324 -1173
rect 290 -1275 324 -1241
rect 290 -1343 324 -1309
rect 290 -1411 324 -1377
rect 290 -1479 324 -1445
rect 290 -1547 324 -1513
rect -221 -1662 -187 -1628
rect -153 -1662 -119 -1628
rect -85 -1662 -51 -1628
rect -17 -1662 17 -1628
rect 51 -1662 85 -1628
rect 119 -1662 153 -1628
rect 187 -1662 221 -1628
<< xpolycontact >>
rect -194 1100 -124 1532
rect -194 -1532 -124 -1100
rect 124 1100 194 1532
rect 124 -1532 194 -1100
<< xpolyres >>
rect -194 -1100 -124 1100
rect 124 -1100 194 1100
<< locali >>
rect -324 1628 -221 1662
rect -187 1628 -153 1662
rect -119 1628 -85 1662
rect -51 1628 -17 1662
rect 17 1628 51 1662
rect 85 1628 119 1662
rect 153 1628 187 1662
rect 221 1628 324 1662
rect -324 1547 -290 1628
rect 290 1547 324 1628
rect -324 1479 -290 1513
rect -324 1411 -290 1445
rect -324 1343 -290 1377
rect -324 1275 -290 1309
rect -324 1207 -290 1241
rect -324 1139 -290 1173
rect -324 1071 -290 1105
rect 290 1479 324 1513
rect 290 1411 324 1445
rect 290 1343 324 1377
rect 290 1275 324 1309
rect 290 1207 324 1241
rect 290 1139 324 1173
rect -324 1003 -290 1037
rect -324 935 -290 969
rect -324 867 -290 901
rect -324 799 -290 833
rect -324 731 -290 765
rect -324 663 -290 697
rect -324 595 -290 629
rect -324 527 -290 561
rect -324 459 -290 493
rect -324 391 -290 425
rect -324 323 -290 357
rect -324 255 -290 289
rect -324 187 -290 221
rect -324 119 -290 153
rect -324 51 -290 85
rect -324 -17 -290 17
rect -324 -85 -290 -51
rect -324 -153 -290 -119
rect -324 -221 -290 -187
rect -324 -289 -290 -255
rect -324 -357 -290 -323
rect -324 -425 -290 -391
rect -324 -493 -290 -459
rect -324 -561 -290 -527
rect -324 -629 -290 -595
rect -324 -697 -290 -663
rect -324 -765 -290 -731
rect -324 -833 -290 -799
rect -324 -901 -290 -867
rect -324 -969 -290 -935
rect -324 -1037 -290 -1003
rect -324 -1105 -290 -1071
rect 290 1071 324 1105
rect 290 1003 324 1037
rect 290 935 324 969
rect 290 867 324 901
rect 290 799 324 833
rect 290 731 324 765
rect 290 663 324 697
rect 290 595 324 629
rect 290 527 324 561
rect 290 459 324 493
rect 290 391 324 425
rect 290 323 324 357
rect 290 255 324 289
rect 290 187 324 221
rect 290 119 324 153
rect 290 51 324 85
rect 290 -17 324 17
rect 290 -85 324 -51
rect 290 -153 324 -119
rect 290 -221 324 -187
rect 290 -289 324 -255
rect 290 -357 324 -323
rect 290 -425 324 -391
rect 290 -493 324 -459
rect 290 -561 324 -527
rect 290 -629 324 -595
rect 290 -697 324 -663
rect 290 -765 324 -731
rect 290 -833 324 -799
rect 290 -901 324 -867
rect 290 -969 324 -935
rect 290 -1037 324 -1003
rect -324 -1173 -290 -1139
rect -324 -1241 -290 -1207
rect -324 -1309 -290 -1275
rect -324 -1377 -290 -1343
rect -324 -1445 -290 -1411
rect -324 -1513 -290 -1479
rect 290 -1105 324 -1071
rect 290 -1173 324 -1139
rect 290 -1241 324 -1207
rect 290 -1309 324 -1275
rect 290 -1377 324 -1343
rect 290 -1445 324 -1411
rect 290 -1513 324 -1479
rect -324 -1628 -290 -1547
rect 290 -1628 324 -1547
rect -324 -1662 -221 -1628
rect -187 -1662 -153 -1628
rect -119 -1662 -85 -1628
rect -51 -1662 -17 -1628
rect 17 -1662 51 -1628
rect 85 -1662 119 -1628
rect 153 -1662 187 -1628
rect 221 -1662 324 -1628
<< properties >>
string FIXED_BBOX -306 -1644 306 1644
<< end >>
