magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< nwell >>
rect 5184 2660 5398 2676
rect -152 2404 5398 2660
rect -152 2384 5370 2404
<< nsubdiff >>
rect -84 2547 5344 2612
rect -84 2513 209 2547
rect 243 2543 1223 2547
rect 243 2513 517 2543
rect -84 2509 517 2513
rect 551 2509 859 2543
rect 893 2513 1223 2543
rect 1257 2543 1953 2547
rect 1257 2513 1575 2543
rect 893 2509 1575 2513
rect 1609 2513 1953 2543
rect 1987 2543 2647 2547
rect 1987 2513 2273 2543
rect 1609 2509 2273 2513
rect 2307 2513 2647 2543
rect 2681 2513 2993 2547
rect 3027 2543 4861 2547
rect 3027 2537 4371 2543
rect 3027 2513 3709 2537
rect 2307 2509 3709 2513
rect -84 2503 3709 2509
rect 3743 2509 4371 2537
rect 4405 2513 4861 2543
rect 4895 2513 5344 2547
rect 4405 2509 5344 2513
rect 3743 2503 5344 2509
rect -84 2452 5344 2503
<< nsubdiffcont >>
rect 209 2513 243 2547
rect 517 2509 551 2543
rect 859 2509 893 2543
rect 1223 2513 1257 2547
rect 1575 2509 1609 2543
rect 1953 2513 1987 2547
rect 2273 2509 2307 2543
rect 2647 2513 2681 2547
rect 2993 2513 3027 2547
rect 3709 2503 3743 2537
rect 4371 2509 4405 2543
rect 4861 2513 4895 2547
<< locali >>
rect 3882 2576 3966 2580
rect -20 2560 5316 2576
rect -20 2554 3907 2560
rect -20 2550 1771 2554
rect -20 2547 369 2550
rect -20 2544 209 2547
rect -20 2510 81 2544
rect 115 2513 209 2544
rect 243 2516 369 2547
rect 403 2543 693 2550
rect 403 2516 517 2543
rect 243 2513 517 2516
rect 115 2510 517 2513
rect -20 2509 517 2510
rect 551 2516 693 2543
rect 727 2543 1041 2550
rect 727 2516 859 2543
rect 551 2509 859 2516
rect 893 2516 1041 2543
rect 1075 2547 1415 2550
rect 1075 2516 1223 2547
rect 893 2513 1223 2516
rect 1257 2516 1415 2547
rect 1449 2543 1771 2550
rect 1449 2516 1575 2543
rect 1257 2513 1575 2516
rect 893 2509 1575 2513
rect 1609 2520 1771 2543
rect 1805 2550 2829 2554
rect 1805 2547 2509 2550
rect 1805 2520 1953 2547
rect 1609 2513 1953 2520
rect 1987 2544 2509 2547
rect 1987 2513 2087 2544
rect 1609 2510 2087 2513
rect 2121 2543 2509 2544
rect 2121 2510 2273 2543
rect 1609 2509 2273 2510
rect 2307 2516 2509 2543
rect 2543 2547 2829 2550
rect 2543 2516 2647 2547
rect 2307 2513 2647 2516
rect 2681 2520 2829 2547
rect 2863 2550 3907 2554
rect 2863 2547 3143 2550
rect 2863 2520 2993 2547
rect 2681 2513 2993 2520
rect 3027 2516 3143 2547
rect 3177 2516 3495 2550
rect 3529 2537 3907 2550
rect 3529 2516 3709 2537
rect 3027 2513 3709 2516
rect 2307 2509 3709 2513
rect -20 2503 3709 2509
rect 3743 2526 3907 2537
rect 3941 2554 5316 2560
rect 3941 2550 4745 2554
rect 3941 2526 4237 2550
rect 3743 2516 4237 2526
rect 4271 2543 4477 2550
rect 4271 2516 4371 2543
rect 3743 2509 4371 2516
rect 4405 2516 4477 2543
rect 4511 2520 4745 2550
rect 4779 2550 5316 2554
rect 4779 2547 4969 2550
rect 4779 2520 4861 2547
rect 4511 2516 4861 2520
rect 4405 2513 4861 2516
rect 4895 2516 4969 2547
rect 5003 2516 5316 2550
rect 4895 2513 5316 2516
rect 4405 2509 5316 2513
rect 3743 2503 5316 2509
rect -20 2474 5316 2503
rect -8 2339 5311 2474
rect 1204 2314 1264 2339
rect 159 2213 176 2247
rect 210 2213 227 2247
rect 317 2213 334 2247
rect 368 2213 385 2247
rect 475 2213 492 2247
rect 526 2213 543 2247
rect 633 2213 650 2247
rect 684 2213 701 2247
rect 791 2213 808 2247
rect 842 2213 859 2247
rect 949 2213 966 2247
rect 1000 2213 1017 2247
rect 1107 2213 1124 2247
rect 1158 2213 1175 2247
rect 1265 2213 1282 2247
rect 1316 2213 1333 2247
rect 1423 2213 1440 2247
rect 1474 2213 1491 2247
rect 1581 2213 1598 2247
rect 1632 2213 1649 2247
rect 1739 2213 1756 2247
rect 1790 2213 1807 2247
rect 1897 2213 1914 2247
rect 1948 2213 1965 2247
rect 2055 2213 2072 2247
rect 2106 2213 2123 2247
rect 2213 2213 2230 2247
rect 2264 2213 2281 2247
rect 2371 2213 2388 2247
rect 2422 2213 2439 2247
rect 98 2052 136 2070
rect 98 2018 100 2052
rect 134 2018 136 2052
rect 98 2000 136 2018
rect 414 2060 452 2078
rect 414 2026 416 2060
rect 450 2026 452 2060
rect 414 2008 452 2026
rect 726 2060 764 2078
rect 726 2026 728 2060
rect 762 2026 764 2060
rect 726 2008 764 2026
rect 1044 2066 1082 2084
rect 1044 2032 1046 2066
rect 1080 2032 1082 2066
rect 1044 2014 1082 2032
rect 1358 2058 1396 2076
rect 1358 2024 1360 2058
rect 1394 2024 1396 2058
rect 1358 2006 1396 2024
rect 1676 2054 1714 2072
rect 1676 2020 1678 2054
rect 1712 2020 1714 2054
rect 1676 2002 1714 2020
rect 1992 2060 2030 2078
rect 1992 2026 1994 2060
rect 2028 2026 2030 2060
rect 1992 2008 2030 2026
rect 2308 2064 2346 2082
rect 2308 2030 2310 2064
rect 2344 2030 2346 2064
rect 2308 2012 2346 2030
rect 252 1798 290 1816
rect 252 1764 254 1798
rect 288 1764 290 1798
rect 252 1746 290 1764
rect 566 1802 604 1820
rect 566 1768 568 1802
rect 602 1768 604 1802
rect 566 1750 604 1768
rect 888 1800 926 1818
rect 888 1766 890 1800
rect 924 1766 926 1800
rect 888 1748 926 1766
rect 1204 1804 1242 1822
rect 1204 1770 1206 1804
rect 1240 1770 1242 1804
rect 1204 1752 1242 1770
rect 1522 1808 1560 1826
rect 1522 1774 1524 1808
rect 1558 1774 1560 1808
rect 1522 1756 1560 1774
rect 1834 1808 1872 1826
rect 1834 1774 1836 1808
rect 1870 1774 1872 1808
rect 1834 1756 1872 1774
rect 2156 1808 2194 1826
rect 2156 1774 2158 1808
rect 2192 1774 2194 1808
rect 2156 1756 2194 1774
rect 2466 1804 2504 1822
rect 2466 1770 2468 1804
rect 2502 1770 2504 1804
rect 2466 1752 2504 1770
rect 2371 85 2388 119
rect 2422 85 2439 119
rect 2584 -16 2703 2339
rect 3746 2322 3806 2339
rect 2860 2218 2877 2252
rect 2911 2218 2928 2252
rect 3018 2218 3035 2252
rect 3069 2218 3086 2252
rect 3176 2218 3193 2252
rect 3227 2218 3244 2252
rect 3334 2218 3351 2252
rect 3385 2218 3402 2252
rect 3492 2218 3509 2252
rect 3543 2218 3560 2252
rect 3650 2218 3667 2252
rect 3701 2218 3718 2252
rect 3808 2218 3825 2252
rect 3859 2218 3876 2252
rect 3966 2218 3983 2252
rect 4017 2218 4034 2252
rect 4124 2218 4141 2252
rect 4175 2218 4192 2252
rect 4282 2218 4299 2252
rect 4333 2218 4350 2252
rect 4440 2218 4457 2252
rect 4491 2218 4508 2252
rect 4598 2218 4615 2252
rect 4649 2218 4666 2252
rect 4756 2218 4773 2252
rect 4807 2218 4824 2252
rect 4914 2218 4931 2252
rect 4965 2218 4982 2252
rect 5072 2218 5089 2252
rect 5123 2218 5140 2252
rect 2796 2026 2832 2060
rect 2796 1992 2797 2026
rect 2831 1992 2832 2026
rect 2796 1958 2832 1992
rect 3110 2040 3146 2074
rect 3110 2006 3111 2040
rect 3145 2006 3146 2040
rect 3110 1972 3146 2006
rect 3270 2004 3304 2088
rect 3428 2040 3464 2074
rect 3428 2006 3429 2040
rect 3463 2006 3464 2040
rect 3586 2012 3620 2096
rect 3746 2036 3782 2070
rect 3428 1972 3464 2006
rect 3746 2002 3747 2036
rect 3781 2002 3782 2036
rect 3902 2016 3936 2100
rect 4058 2042 4094 2076
rect 3746 1968 3782 2002
rect 4058 2008 4059 2042
rect 4093 2008 4094 2042
rect 4058 1974 4094 2008
rect 4374 2044 4410 2078
rect 4374 2010 4375 2044
rect 4409 2010 4410 2044
rect 4374 1976 4410 2010
rect 4690 2036 4726 2070
rect 4690 2002 4691 2036
rect 4725 2002 4726 2036
rect 4690 1968 4726 2002
rect 5012 2040 5048 2074
rect 5012 2006 5013 2040
rect 5047 2006 5048 2040
rect 5012 1972 5048 2006
rect 3268 1857 3302 1858
rect 2956 1849 2990 1850
rect 2956 1777 2990 1815
rect 3902 1855 3936 1856
rect 3268 1785 3302 1823
rect 3268 1750 3302 1751
rect 3586 1853 3620 1854
rect 3586 1781 3620 1819
rect 3902 1783 3936 1821
rect 3902 1748 3936 1749
rect 4222 1855 4256 1856
rect 4222 1783 4256 1821
rect 4222 1748 4256 1749
rect 4536 1849 4570 1850
rect 4536 1777 4570 1815
rect 3586 1746 3620 1747
rect 2956 1742 2990 1743
rect 4536 1742 4570 1743
rect 4852 1849 4886 1850
rect 4852 1777 4886 1815
rect 4852 1742 4886 1743
rect 5168 1849 5202 1850
rect 5168 1777 5202 1815
rect 5168 1742 5202 1743
rect 2392 -402 2405 -368
rect 2439 -402 2452 -368
rect 2894 -404 2907 -370
rect 2941 -404 2954 -370
rect 2392 -490 2405 -456
rect 2439 -490 2452 -456
rect 2894 -492 2907 -458
rect 2941 -492 2954 -458
rect 2396 -602 2412 -568
rect 2446 -602 2462 -568
rect 2892 -606 2908 -572
rect 2942 -606 2958 -572
rect 2642 -1016 2648 -982
rect 2682 -1016 2688 -982
rect 1478 -1586 1487 -1552
rect 1521 -1586 1530 -1552
rect 1810 -1592 1819 -1558
rect 1853 -1592 1862 -1558
rect 2292 -1592 2301 -1558
rect 2335 -1592 2344 -1558
rect 2944 -1586 2953 -1552
rect 2987 -1586 2996 -1552
rect 3530 -1590 3539 -1556
rect 3573 -1590 3582 -1556
rect 3848 -1588 3857 -1554
rect 3891 -1588 3900 -1554
<< viali >>
rect 81 2510 115 2544
rect 369 2516 403 2550
rect 693 2516 727 2550
rect 1041 2516 1075 2550
rect 1415 2516 1449 2550
rect 1771 2520 1805 2554
rect 2087 2510 2121 2544
rect 2509 2516 2543 2550
rect 2829 2520 2863 2554
rect 3143 2516 3177 2550
rect 3495 2516 3529 2550
rect 3907 2526 3941 2560
rect 4237 2516 4271 2550
rect 4477 2516 4511 2550
rect 4745 2520 4779 2554
rect 4969 2516 5003 2550
rect 176 2213 210 2247
rect 334 2213 368 2247
rect 492 2213 526 2247
rect 650 2213 684 2247
rect 808 2213 842 2247
rect 966 2213 1000 2247
rect 1124 2213 1158 2247
rect 1282 2213 1316 2247
rect 1440 2213 1474 2247
rect 1598 2213 1632 2247
rect 1756 2213 1790 2247
rect 1914 2213 1948 2247
rect 2072 2213 2106 2247
rect 2230 2213 2264 2247
rect 2388 2213 2422 2247
rect 100 2018 134 2052
rect 416 2026 450 2060
rect 728 2026 762 2060
rect 1046 2032 1080 2066
rect 1360 2024 1394 2058
rect 1678 2020 1712 2054
rect 1994 2026 2028 2060
rect 2310 2030 2344 2064
rect 254 1764 288 1798
rect 568 1768 602 1802
rect 890 1766 924 1800
rect 1206 1770 1240 1804
rect 1524 1774 1558 1808
rect 1836 1774 1870 1808
rect 2158 1774 2192 1808
rect 2468 1770 2502 1804
rect 176 85 210 119
rect 334 85 368 119
rect 492 85 526 119
rect 650 85 684 119
rect 808 85 842 119
rect 966 85 1000 119
rect 1124 85 1158 119
rect 1282 85 1316 119
rect 1440 85 1474 119
rect 1598 85 1632 119
rect 1756 85 1790 119
rect 1914 85 1948 119
rect 2072 85 2106 119
rect 2230 85 2264 119
rect 2388 85 2422 119
rect 2877 2218 2911 2252
rect 3035 2218 3069 2252
rect 3193 2218 3227 2252
rect 3351 2218 3385 2252
rect 3509 2218 3543 2252
rect 3667 2218 3701 2252
rect 3825 2218 3859 2252
rect 3983 2218 4017 2252
rect 4141 2218 4175 2252
rect 4299 2218 4333 2252
rect 4457 2218 4491 2252
rect 4615 2218 4649 2252
rect 4773 2218 4807 2252
rect 4931 2218 4965 2252
rect 5089 2218 5123 2252
rect 2797 1992 2831 2026
rect 3111 2006 3145 2040
rect 3429 2006 3463 2040
rect 3747 2002 3781 2036
rect 4059 2008 4093 2042
rect 4375 2010 4409 2044
rect 4691 2002 4725 2036
rect 5013 2006 5047 2040
rect 2956 1815 2990 1849
rect 2956 1743 2990 1777
rect 3268 1823 3302 1857
rect 3268 1751 3302 1785
rect 3586 1819 3620 1853
rect 3586 1747 3620 1781
rect 3902 1821 3936 1855
rect 3902 1749 3936 1783
rect 4222 1821 4256 1855
rect 4222 1749 4256 1783
rect 4536 1815 4570 1849
rect 4536 1743 4570 1777
rect 4852 1815 4886 1849
rect 4852 1743 4886 1777
rect 5168 1815 5202 1849
rect 5168 1743 5202 1777
rect 2929 90 2963 124
rect 3035 90 3069 124
rect 3193 90 3227 124
rect 3351 90 3385 124
rect 3509 90 3543 124
rect 3667 90 3701 124
rect 3825 90 3859 124
rect 3983 90 4017 124
rect 4141 90 4175 124
rect 4299 90 4333 124
rect 4457 90 4491 124
rect 4615 90 4649 124
rect 4773 90 4807 124
rect 4931 90 4965 124
rect 5089 90 5123 124
rect 2405 -402 2439 -368
rect 2907 -404 2941 -370
rect 2405 -490 2439 -456
rect 2907 -492 2941 -458
rect 2412 -602 2446 -568
rect 2908 -606 2942 -572
rect 2648 -1016 2682 -982
rect 1487 -1586 1521 -1552
rect 1819 -1592 1853 -1558
rect 2301 -1592 2335 -1558
rect 2953 -1586 2987 -1552
rect 3539 -1590 3573 -1556
rect 3857 -1588 3891 -1554
<< metal1 >>
rect -110 2583 5338 2628
rect -110 2544 93 2583
rect 145 2560 5338 2583
rect 145 2554 3907 2560
rect 145 2550 1771 2554
rect -110 2510 81 2544
rect 145 2531 369 2550
rect 115 2519 369 2531
rect 145 2516 369 2519
rect 403 2516 693 2550
rect 727 2516 1041 2550
rect 1075 2516 1415 2550
rect 1449 2520 1771 2550
rect 1805 2550 2829 2554
rect 1805 2544 2509 2550
rect 1805 2520 2087 2544
rect 1449 2516 2087 2520
rect 145 2510 2087 2516
rect 2121 2516 2509 2544
rect 2543 2520 2829 2550
rect 2863 2550 3907 2554
rect 2863 2520 3143 2550
rect 2543 2516 3143 2520
rect 3177 2516 3495 2550
rect 3529 2526 3907 2550
rect 3941 2554 5338 2560
rect 3941 2550 4745 2554
rect 3941 2526 4237 2550
rect 3529 2516 4237 2526
rect 4271 2516 4477 2550
rect 4511 2520 4745 2550
rect 4779 2550 5338 2554
rect 4779 2520 4969 2550
rect 4511 2516 4969 2520
rect 5003 2546 5338 2550
rect 5003 2516 5157 2546
rect 2121 2510 5157 2516
rect -110 2467 93 2510
rect 145 2494 5157 2510
rect 5209 2494 5338 2546
rect 145 2467 5338 2494
rect -110 2436 5338 2467
rect 2830 2274 5170 2278
rect 132 2252 5170 2274
rect 132 2247 2877 2252
rect 132 2213 176 2247
rect 210 2213 334 2247
rect 368 2213 492 2247
rect 526 2213 650 2247
rect 684 2213 808 2247
rect 842 2213 966 2247
rect 1000 2213 1124 2247
rect 1158 2213 1282 2247
rect 1316 2213 1440 2247
rect 1474 2213 1598 2247
rect 1632 2213 1756 2247
rect 1790 2213 1914 2247
rect 1948 2213 2072 2247
rect 2106 2213 2230 2247
rect 2264 2213 2388 2247
rect 2422 2218 2877 2247
rect 2911 2218 3035 2252
rect 3069 2218 3193 2252
rect 3227 2218 3351 2252
rect 3385 2218 3509 2252
rect 3543 2218 3667 2252
rect 3701 2218 3825 2252
rect 3859 2218 3983 2252
rect 4017 2218 4141 2252
rect 4175 2218 4299 2252
rect 4333 2218 4457 2252
rect 4491 2218 4615 2252
rect 4649 2218 4773 2252
rect 4807 2218 4931 2252
rect 4965 2218 5089 2252
rect 5123 2218 5170 2252
rect 2422 2213 5170 2218
rect 132 2200 5170 2213
rect 2350 2196 3320 2200
rect 26 2110 234 2124
rect 26 2103 2356 2110
rect 26 2051 93 2103
rect 145 2066 2356 2103
rect 145 2060 1046 2066
rect 145 2051 416 2060
rect 26 2039 100 2051
rect 134 2039 416 2051
rect 26 1987 93 2039
rect 145 2026 416 2039
rect 450 2026 728 2060
rect 762 2032 1046 2060
rect 1080 2064 2356 2066
rect 1080 2060 2310 2064
rect 1080 2058 1994 2060
rect 1080 2032 1360 2058
rect 762 2026 1360 2032
rect 145 2024 1360 2026
rect 1394 2054 1994 2058
rect 1394 2024 1678 2054
rect 145 2020 1678 2024
rect 1712 2026 1994 2054
rect 2028 2030 2310 2060
rect 2344 2030 2356 2064
rect 2028 2026 2356 2030
rect 1712 2020 2356 2026
rect 145 1987 2356 2020
rect 26 1962 2356 1987
rect 26 1944 234 1962
rect 2750 2084 2874 2086
rect 2750 2044 5062 2084
rect 2750 2042 4375 2044
rect 2750 2040 4059 2042
rect 2750 2026 3111 2040
rect 2750 1992 2797 2026
rect 2831 2006 3111 2026
rect 3145 2006 3429 2040
rect 3463 2036 4059 2040
rect 3463 2006 3747 2036
rect 2831 2002 3747 2006
rect 3781 2008 4059 2036
rect 4093 2010 4375 2042
rect 4409 2040 5062 2044
rect 4409 2036 5013 2040
rect 4409 2010 4691 2036
rect 4093 2008 4691 2010
rect 3781 2002 4691 2008
rect 4725 2006 5013 2036
rect 5047 2006 5062 2040
rect 4725 2002 5062 2006
rect 2831 1992 5062 2002
rect 2750 1950 5062 1992
rect 2426 1864 2546 1870
rect 238 1808 2546 1864
rect 2750 1832 2874 1950
rect 5108 1864 5260 1878
rect 238 1804 1524 1808
rect 238 1802 1206 1804
rect 238 1798 568 1802
rect 238 1764 254 1798
rect 288 1768 568 1798
rect 602 1800 1206 1802
rect 602 1768 890 1800
rect 288 1766 890 1768
rect 924 1770 1206 1800
rect 1240 1774 1524 1804
rect 1558 1774 1836 1808
rect 1870 1774 2158 1808
rect 2192 1804 2546 1808
rect 2192 1774 2468 1804
rect 1240 1770 2468 1774
rect 2502 1770 2546 1804
rect 924 1766 2546 1770
rect 288 1764 2546 1766
rect 238 1700 2546 1764
rect 2426 134 2546 1700
rect 2352 129 2546 134
rect 121 124 2546 129
rect 121 69 156 124
rect 2419 119 2546 124
rect 2422 85 2546 119
rect 2419 69 2546 85
rect 121 68 2546 69
rect 2352 64 2546 68
rect 2426 -152 2546 64
rect 2372 -178 2546 -152
rect 2738 62 2874 1832
rect 2944 1857 5260 1864
rect 2944 1849 3268 1857
rect 2944 1815 2956 1849
rect 2990 1823 3268 1849
rect 3302 1855 5260 1857
rect 3302 1853 3902 1855
rect 3302 1823 3586 1853
rect 2990 1819 3586 1823
rect 3620 1821 3902 1853
rect 3936 1821 4222 1855
rect 4256 1849 5260 1855
rect 4256 1821 4536 1849
rect 3620 1819 4536 1821
rect 2990 1815 4536 1819
rect 4570 1815 4852 1849
rect 4886 1815 5168 1849
rect 5202 1820 5260 1849
rect 2944 1785 5175 1815
rect 2944 1777 3268 1785
rect 2944 1743 2956 1777
rect 2990 1751 3268 1777
rect 3302 1783 5175 1785
rect 3302 1781 3902 1783
rect 3302 1751 3586 1781
rect 2990 1747 3586 1751
rect 3620 1749 3902 1781
rect 3936 1749 4222 1783
rect 4256 1777 5175 1783
rect 4256 1749 4536 1777
rect 3620 1747 4536 1749
rect 2990 1743 4536 1747
rect 4570 1743 4852 1777
rect 4886 1743 5168 1777
rect 5227 1768 5260 1820
rect 5202 1743 5260 1768
rect 2944 1734 5260 1743
rect 5108 1724 5260 1734
rect 2916 124 5163 131
rect 2916 90 2929 124
rect 2963 123 3035 124
rect 3069 123 3193 124
rect 3227 123 3351 124
rect 3385 123 3509 124
rect 3543 123 3667 124
rect 3701 123 3825 124
rect 3859 123 3983 124
rect 4017 123 4141 124
rect 4175 123 4299 124
rect 4333 123 4457 124
rect 4491 123 4615 124
rect 4649 123 4773 124
rect 4807 123 4931 124
rect 4965 123 5089 124
rect 5083 90 5089 123
rect 5123 90 5163 124
rect 2916 78 2953 90
rect 2943 70 2953 78
rect 5083 78 5163 90
rect 5083 70 5093 78
rect 2738 -136 2862 62
rect 2372 -352 2474 -178
rect 2738 -192 2976 -136
rect 2846 -196 2976 -192
rect 2372 -368 2478 -352
rect 2372 -402 2405 -368
rect 2439 -402 2478 -368
rect 2372 -406 2478 -402
rect 2378 -410 2478 -406
rect 2874 -370 2976 -196
rect 2874 -404 2907 -370
rect 2941 -404 2976 -370
rect 2874 -410 2976 -404
rect 2366 -456 2476 -450
rect 2366 -490 2405 -456
rect 2439 -490 2476 -456
rect 2366 -558 2476 -490
rect 2872 -458 2982 -452
rect 2872 -492 2907 -458
rect 2941 -492 2982 -458
rect 2872 -558 2982 -492
rect 2362 -568 2982 -558
rect 2362 -602 2412 -568
rect 2446 -572 2982 -568
rect 2446 -602 2908 -572
rect 2362 -606 2908 -602
rect 2942 -606 2982 -572
rect 2362 -620 2982 -606
rect 2622 -728 2708 -620
rect 2622 -982 2706 -728
rect 2622 -1016 2648 -982
rect 2682 -1016 2706 -982
rect 2622 -1018 2706 -1016
rect 2626 -1022 2706 -1018
rect 1170 -1552 4300 -1522
rect 1170 -1586 1487 -1552
rect 1521 -1558 2953 -1552
rect 1521 -1586 1819 -1558
rect 1170 -1592 1819 -1586
rect 1853 -1592 2301 -1558
rect 2335 -1586 2953 -1558
rect 2987 -1554 4300 -1552
rect 2987 -1556 3857 -1554
rect 2987 -1586 3539 -1556
rect 2335 -1590 3539 -1586
rect 3573 -1588 3857 -1556
rect 3891 -1588 4300 -1554
rect 3573 -1590 4300 -1588
rect 2335 -1592 4300 -1590
rect 1170 -1748 4300 -1592
<< rmetal1 >>
rect 234 1960 2356 1962
<< via1 >>
rect 93 2544 145 2583
rect 93 2531 115 2544
rect 115 2531 145 2544
rect 93 2510 115 2519
rect 115 2510 145 2519
rect 93 2467 145 2510
rect 5157 2494 5209 2546
rect 93 2052 145 2103
rect 93 2051 100 2052
rect 100 2051 134 2052
rect 134 2051 145 2052
rect 93 2018 100 2039
rect 100 2018 134 2039
rect 134 2018 145 2039
rect 93 1987 145 2018
rect 156 119 2419 124
rect 156 85 176 119
rect 176 85 210 119
rect 210 85 334 119
rect 334 85 368 119
rect 368 85 492 119
rect 492 85 526 119
rect 526 85 650 119
rect 650 85 684 119
rect 684 85 808 119
rect 808 85 842 119
rect 842 85 966 119
rect 966 85 1000 119
rect 1000 85 1124 119
rect 1124 85 1158 119
rect 1158 85 1282 119
rect 1282 85 1316 119
rect 1316 85 1440 119
rect 1440 85 1474 119
rect 1474 85 1598 119
rect 1598 85 1632 119
rect 1632 85 1756 119
rect 1756 85 1790 119
rect 1790 85 1914 119
rect 1914 85 1948 119
rect 1948 85 2072 119
rect 2072 85 2106 119
rect 2106 85 2230 119
rect 2230 85 2264 119
rect 2264 85 2388 119
rect 2388 85 2419 119
rect 156 69 2419 85
rect 5175 1815 5202 1820
rect 5202 1815 5227 1820
rect 5175 1777 5227 1815
rect 5175 1768 5202 1777
rect 5202 1768 5227 1777
rect 2953 90 2963 123
rect 2963 90 3035 123
rect 3035 90 3069 123
rect 3069 90 3193 123
rect 3193 90 3227 123
rect 3227 90 3351 123
rect 3351 90 3385 123
rect 3385 90 3509 123
rect 3509 90 3543 123
rect 3543 90 3667 123
rect 3667 90 3701 123
rect 3701 90 3825 123
rect 3825 90 3859 123
rect 3859 90 3983 123
rect 3983 90 4017 123
rect 4017 90 4141 123
rect 4141 90 4175 123
rect 4175 90 4299 123
rect 4299 90 4333 123
rect 4333 90 4457 123
rect 4457 90 4491 123
rect 4491 90 4615 123
rect 4615 90 4649 123
rect 4649 90 4773 123
rect 4773 90 4807 123
rect 4807 90 4931 123
rect 4931 90 4965 123
rect 4965 90 5083 123
rect 2953 70 5083 90
<< metal2 >>
rect 44 2583 194 2618
rect 44 2531 93 2583
rect 145 2531 194 2583
rect 44 2519 194 2531
rect 44 2467 93 2519
rect 145 2467 194 2519
rect 44 2103 194 2467
rect 44 2051 93 2103
rect 145 2051 194 2103
rect 44 2039 194 2051
rect 44 1987 93 2039
rect 145 1987 194 2039
rect 44 1938 194 1987
rect 5116 2546 5276 2584
rect 5116 2494 5157 2546
rect 5209 2494 5276 2546
rect 5116 1820 5276 2494
rect 5116 1768 5175 1820
rect 5227 1768 5276 1820
rect 5116 1724 5276 1768
rect 156 131 2419 134
rect 2953 131 5083 133
rect 138 124 5163 131
rect 138 69 156 124
rect 2419 123 5163 124
rect 2419 70 2953 123
rect 5083 70 5163 123
rect 2419 69 5163 70
rect 138 64 5163 69
rect 156 59 2419 64
rect 2953 60 5083 64
use sky130_fd_pr__nfet_01v8_lvt_69NU8X  sky130_fd_pr__nfet_01v8_lvt_69NU8X_0
timestamp 1699818132
transform 0 1 2704 -1 0 -1228
box -360 -1434 360 1434
use sky130_fd_pr__nfet_01v8_lvt_D42ZUM  sky130_fd_pr__nfet_01v8_lvt_D42ZUM_0
timestamp 1699818132
transform 0 1 2924 -1 0 -431
box -175 -216 175 216
use sky130_fd_pr__nfet_01v8_lvt_D42ZUM  sky130_fd_pr__nfet_01v8_lvt_D42ZUM_1
timestamp 1699818132
transform 0 1 2422 -1 0 -429
box -175 -216 175 216
use sky130_fd_pr__pfet_01v8_NC6LGM  sky130_fd_pr__pfet_01v8_NC6LGM_0
timestamp 1699818132
transform 1 0 1299 0 1 1166
box -1352 -1219 1352 1219
use sky130_fd_pr__pfet_01v8_NC6LGM  sky130_fd_pr__pfet_01v8_NC6LGM_1
timestamp 1699818132
transform 1 0 4000 0 1 1171
box -1352 -1219 1352 1219
<< labels >>
rlabel metal1 s 2652 -744 2684 -700 4 Itail_b
rlabel metal1 s 2356 2494 2412 2550 4 Vdd
port 1 nsew
rlabel metal1 s 2460 -134 2516 -78 4 ON2b
port 2 nsew
rlabel metal1 s 2778 -132 2834 -76 4 ON1b
port 3 nsew
rlabel metal1 s 2664 -1694 2750 -1640 4 Gnd
port 4 nsew
<< end >>
