magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< nwell >>
rect 15607 3090 19358 3322
rect 15572 3076 19358 3090
rect 15566 2980 19358 3076
rect 15566 2796 19158 2980
rect 15566 2782 19152 2796
<< psubdiff >>
rect 16126 2266 16150 2382
rect 19262 2266 19286 2382
<< nsubdiff >>
rect 16104 3192 19252 3232
rect 16104 3108 16152 3192
rect 19214 3108 19252 3192
rect 16104 3074 19252 3108
<< psubdiffcont >>
rect 16150 2266 19262 2382
<< nsubdiffcont >>
rect 16152 3108 19214 3192
<< locali >>
rect 16120 3192 19244 3200
rect 43 3079 352 3136
rect 16120 3108 16152 3192
rect 19214 3108 19244 3192
rect 16120 3104 19244 3108
rect 43 2937 64 3079
rect 323 2937 352 3079
rect 43 2884 352 2937
rect 7748 2838 7824 2902
rect 8346 2852 8426 2902
rect 17930 2738 17970 2740
rect 17046 2717 17080 2718
rect 16244 2701 16278 2702
rect 16152 2699 16186 2700
rect 17930 2704 17933 2738
rect 17967 2704 17970 2738
rect 17930 2702 17970 2704
rect 17046 2682 17080 2683
rect 16244 2666 16278 2667
rect 16152 2664 16186 2665
rect 19050 2622 19088 2626
rect 17138 2620 17178 2622
rect 17138 2586 17141 2620
rect 17175 2586 17178 2620
rect 17138 2584 17178 2586
rect 18020 2620 18060 2622
rect 18020 2586 18023 2620
rect 18057 2586 18060 2620
rect 18020 2584 18060 2586
rect 19050 2588 19052 2622
rect 19086 2588 19088 2622
rect 19050 2584 19088 2588
rect 12568 2434 12602 2438
rect 12568 2421 12622 2434
rect 12568 2387 12576 2421
rect 12610 2387 12622 2421
rect 12568 2368 12622 2387
rect 13300 2386 13303 2420
rect 13337 2386 13340 2420
rect 12568 2364 12602 2368
rect 16134 2266 16150 2382
rect 19262 2266 19278 2382
rect 8667 1367 8849 1674
rect 9138 1367 9320 1675
rect 11652 1516 11688 1528
rect 11652 1482 11653 1516
rect 11687 1482 11688 1516
rect 11652 1470 11688 1482
rect 8667 1155 9320 1367
rect 11738 1358 11745 1392
rect 11779 1358 11817 1392
rect 11851 1358 11889 1392
rect 11923 1358 11961 1392
rect 11995 1358 12033 1392
rect 12067 1358 12105 1392
rect 12139 1358 12177 1392
rect 12211 1358 12249 1392
rect 12283 1358 12321 1392
rect 12355 1358 12393 1392
rect 12427 1358 12465 1392
rect 12499 1358 12537 1392
rect 12571 1358 12609 1392
rect 12643 1358 12681 1392
rect 12715 1358 12753 1392
rect 12787 1358 12825 1392
rect 12859 1358 12897 1392
rect 12931 1358 12969 1392
rect 13003 1358 13041 1392
rect 13075 1358 13113 1392
rect 13147 1358 13185 1392
rect 13219 1358 13257 1392
rect 13291 1358 13329 1392
rect 13363 1358 13401 1392
rect 13435 1358 13473 1392
rect 13507 1358 13545 1392
rect 13579 1358 13617 1392
rect 13651 1358 13689 1392
rect 13723 1358 13761 1392
rect 13795 1358 13833 1392
rect 13867 1358 13905 1392
rect 13939 1358 13977 1392
rect 14011 1358 14049 1392
rect 14083 1358 14121 1392
rect 14155 1358 14193 1392
rect 14227 1358 14234 1392
rect 8667 954 8683 1155
rect 9300 954 9320 1155
rect 8667 939 9320 954
rect 8667 937 8849 939
rect 9138 938 9320 939
rect 5302 78 5333 112
rect 5367 78 5405 112
rect 5439 78 5477 112
rect 5511 78 5549 112
rect 5583 78 5621 112
rect 5655 78 5693 112
rect 5727 78 5758 112
rect 2438 24 2469 58
rect 2503 24 2541 58
rect 2575 24 2613 58
rect 2647 24 2685 58
rect 2719 24 2757 58
rect 2791 24 2829 58
rect 2863 24 2894 58
<< viali >>
rect 16152 3108 19214 3192
rect 64 2937 323 3079
rect 16152 2665 16186 2699
rect 16244 2667 16278 2701
rect 17046 2683 17080 2717
rect 17933 2704 17967 2738
rect 18956 2714 18990 2748
rect 17141 2586 17175 2620
rect 18023 2586 18057 2620
rect 19052 2588 19086 2622
rect 12576 2387 12610 2421
rect 13303 2386 13337 2420
rect 16150 2266 19262 2382
rect 11653 1482 11687 1516
rect 11745 1358 11779 1392
rect 11817 1358 11851 1392
rect 11889 1358 11923 1392
rect 11961 1358 11995 1392
rect 12033 1358 12067 1392
rect 12105 1358 12139 1392
rect 12177 1358 12211 1392
rect 12249 1358 12283 1392
rect 12321 1358 12355 1392
rect 12393 1358 12427 1392
rect 12465 1358 12499 1392
rect 12537 1358 12571 1392
rect 12609 1358 12643 1392
rect 12681 1358 12715 1392
rect 12753 1358 12787 1392
rect 12825 1358 12859 1392
rect 12897 1358 12931 1392
rect 12969 1358 13003 1392
rect 13041 1358 13075 1392
rect 13113 1358 13147 1392
rect 13185 1358 13219 1392
rect 13257 1358 13291 1392
rect 13329 1358 13363 1392
rect 13401 1358 13435 1392
rect 13473 1358 13507 1392
rect 13545 1358 13579 1392
rect 13617 1358 13651 1392
rect 13689 1358 13723 1392
rect 13761 1358 13795 1392
rect 13833 1358 13867 1392
rect 13905 1358 13939 1392
rect 13977 1358 14011 1392
rect 14049 1358 14083 1392
rect 14121 1358 14155 1392
rect 14193 1358 14227 1392
rect 8683 954 9300 1155
rect 5333 78 5367 112
rect 5405 78 5439 112
rect 5477 78 5511 112
rect 5549 78 5583 112
rect 5621 78 5655 112
rect 5693 78 5727 112
rect 2469 24 2503 58
rect 2541 24 2575 58
rect 2613 24 2647 58
rect 2685 24 2719 58
rect 2757 24 2791 58
rect 2829 24 2863 58
<< metal1 >>
rect 3372 5570 19328 5860
rect 4688 5510 19328 5570
rect 6474 5414 19328 5510
rect 6555 5316 19328 5414
rect 6555 5268 9736 5316
rect 9640 5260 9736 5268
rect 9808 5268 19328 5316
rect 9808 5260 10306 5268
rect 8434 4790 8518 4814
rect 8434 4738 8450 4790
rect 8502 4738 8518 4790
rect 8434 4714 8518 4738
rect 9952 4800 10062 4838
rect 9952 4748 9984 4800
rect 10036 4748 10062 4800
rect 7746 4664 7840 4668
rect 7746 4612 7767 4664
rect 7819 4612 7840 4664
rect 7746 4600 7840 4612
rect 7746 4548 7767 4600
rect 7819 4548 7840 4600
rect 7746 4544 7840 4548
rect 9952 4252 10062 4748
rect 12002 4252 12100 4260
rect 9952 4168 12104 4252
rect 9958 4162 12104 4168
rect 145 3568 257 3582
rect 145 3482 158 3568
rect 244 3482 257 3568
rect 145 3469 257 3482
rect 158 3231 244 3469
rect 52 3079 335 3085
rect 52 2937 64 3079
rect 323 2937 335 3079
rect 8250 3022 8310 3036
rect 7600 3011 7652 3016
rect 7600 2954 7652 2959
rect 8250 2970 8254 3022
rect 8306 2970 8310 3022
rect 8250 2956 8310 2970
rect 8614 3015 8666 3030
rect 8614 2948 8666 2963
rect 52 2931 335 2937
rect 7758 2902 7820 2904
rect 7748 2894 7824 2902
rect 7424 2888 7828 2894
rect 7424 2836 7439 2888
rect 7491 2836 7828 2888
rect 7424 2830 7828 2836
rect 8346 2892 8422 2900
rect 8346 2858 8370 2892
rect 8404 2858 8422 2892
rect 159 2552 245 2790
rect 7390 2726 7484 2730
rect 7390 2674 7414 2726
rect 7466 2714 7484 2726
rect 8346 2714 8422 2858
rect 12002 2780 12100 4162
rect 16062 3192 19328 5268
rect 16062 3108 16152 3192
rect 19214 3108 19328 3192
rect 16062 3017 19328 3108
rect 16062 2940 16236 3017
rect 16332 2936 16982 3017
rect 17212 2996 19270 3017
rect 17212 2992 19176 2996
rect 7466 2674 8424 2714
rect 7390 2672 8424 2674
rect 7390 2656 7484 2672
rect 147 2539 259 2552
rect 147 2453 159 2539
rect 245 2453 259 2539
rect 147 2439 259 2453
rect 9710 2356 9720 2712
rect 9894 2436 9904 2712
rect 12002 2701 12138 2780
rect 18018 2750 19002 2762
rect 17956 2748 19002 2750
rect 17134 2738 18956 2748
rect 17134 2730 17933 2738
rect 16230 2717 17933 2730
rect 12002 2649 12043 2701
rect 12095 2649 12138 2701
rect 12002 2640 12138 2649
rect 13112 2708 15704 2710
rect 13112 2699 16200 2708
rect 13112 2665 16152 2699
rect 16186 2665 16200 2699
rect 13112 2644 16200 2665
rect 16230 2701 17046 2717
rect 16230 2667 16244 2701
rect 16278 2683 17046 2701
rect 17080 2704 17933 2717
rect 17967 2714 18956 2738
rect 18990 2714 19002 2748
rect 17967 2704 19002 2714
rect 17080 2694 19002 2704
rect 17080 2683 18118 2694
rect 16278 2682 18118 2683
rect 16278 2676 17986 2682
rect 16278 2667 17348 2676
rect 16230 2666 17348 2667
rect 16230 2658 17102 2666
rect 12008 2614 12138 2640
rect 19146 2638 19328 2646
rect 18014 2632 19328 2638
rect 17118 2622 19328 2632
rect 17118 2620 19052 2622
rect 17118 2586 17141 2620
rect 17175 2601 18023 2620
rect 17175 2586 17784 2601
rect 17118 2570 17784 2586
rect 17858 2586 18023 2601
rect 18057 2605 19052 2620
rect 18057 2586 18133 2605
rect 17858 2574 18133 2586
rect 18207 2588 19052 2605
rect 19086 2588 19328 2622
rect 18207 2574 19328 2588
rect 17858 2570 18064 2574
rect 19148 2506 19258 2534
rect 16338 2473 16988 2506
rect 17200 2473 19258 2506
rect 12296 2436 12618 2440
rect 13484 2436 13594 2438
rect 9894 2421 12618 2436
rect 9894 2387 12576 2421
rect 12610 2387 12618 2421
rect 9894 2366 12618 2387
rect 13294 2420 13594 2436
rect 16162 2424 19328 2473
rect 13294 2386 13303 2420
rect 13337 2386 13594 2420
rect 13294 2366 13594 2386
rect 9894 2364 12310 2366
rect 9894 2356 9904 2364
rect 4982 1946 5086 2340
rect 8084 2134 8196 2164
rect 8084 2082 8114 2134
rect 8166 2082 8196 2134
rect 8084 2052 8196 2082
rect 13484 2113 13594 2366
rect 13484 2061 13508 2113
rect 13560 2061 13594 2113
rect 13484 2030 13594 2061
rect 16080 2382 19328 2424
rect 16080 2266 16150 2382
rect 19262 2266 19328 2382
rect 4982 1776 7978 1946
rect 9508 1871 9594 1884
rect 9508 1819 9525 1871
rect 9577 1819 9594 1871
rect 9508 1806 9594 1819
rect 5912 1171 7978 1776
rect 8060 1454 8070 1640
rect 8516 1554 8526 1640
rect 8516 1516 11712 1554
rect 8516 1482 11653 1516
rect 11687 1482 11712 1516
rect 8516 1462 11712 1482
rect 8516 1454 8526 1462
rect 11722 1392 14248 1404
rect 11722 1358 11745 1392
rect 11779 1358 11817 1392
rect 11851 1358 11889 1392
rect 11923 1358 11961 1392
rect 11995 1358 12033 1392
rect 12067 1358 12105 1392
rect 12139 1358 12177 1392
rect 12211 1358 12249 1392
rect 12283 1358 12321 1392
rect 12355 1358 12393 1392
rect 12427 1358 12465 1392
rect 12499 1358 12537 1392
rect 12571 1358 12609 1392
rect 12643 1358 12681 1392
rect 12715 1358 12753 1392
rect 12787 1358 12825 1392
rect 12859 1358 12897 1392
rect 12931 1358 12969 1392
rect 13003 1358 13041 1392
rect 13075 1358 13113 1392
rect 13147 1358 13185 1392
rect 13219 1358 13257 1392
rect 13291 1358 13329 1392
rect 13363 1358 13401 1392
rect 13435 1358 13473 1392
rect 13507 1358 13545 1392
rect 13579 1358 13617 1392
rect 13651 1358 13689 1392
rect 13723 1358 13761 1392
rect 13795 1358 13833 1392
rect 13867 1358 13905 1392
rect 13939 1358 13977 1392
rect 14011 1358 14049 1392
rect 14083 1358 14121 1392
rect 14155 1358 14193 1392
rect 14227 1358 14248 1392
rect 11722 1280 14248 1358
rect 16080 1310 19328 2266
rect 11482 1239 11568 1252
rect 14572 1248 19328 1310
rect 11482 1187 11499 1239
rect 11551 1187 11568 1239
rect 11482 1174 11568 1187
rect 14561 1171 19328 1248
rect 5912 1155 19328 1171
rect 5912 954 8683 1155
rect 9300 954 19328 1155
rect 5272 112 5798 123
rect 5272 82 5333 112
rect 2306 78 5333 82
rect 5367 78 5405 112
rect 5439 78 5477 112
rect 5511 78 5549 112
rect 5583 78 5621 112
rect 5655 78 5693 112
rect 5727 82 5798 112
rect 5912 82 19328 954
rect 5727 78 19328 82
rect 2306 58 19328 78
rect 2306 24 2469 58
rect 2503 24 2541 58
rect 2575 24 2613 58
rect 2647 24 2685 58
rect 2719 24 2757 58
rect 2791 24 2829 58
rect 2863 24 19328 58
rect 2306 4 19328 24
<< via1 >>
rect 8450 4738 8502 4790
rect 9984 4748 10036 4800
rect 7767 4612 7819 4664
rect 7767 4548 7819 4600
rect 158 3482 244 3568
rect 64 2937 323 3079
rect 7600 2959 7652 3011
rect 8254 2970 8306 3022
rect 8614 2963 8666 3015
rect 7439 2836 7491 2888
rect 7414 2674 7466 2726
rect 159 2453 245 2539
rect 9720 2356 9894 2712
rect 12043 2649 12095 2701
rect 8114 2082 8166 2134
rect 13508 2061 13560 2113
rect 9525 1819 9577 1871
rect 8070 1454 8516 1640
rect 11499 1187 11551 1239
<< metal2 >>
rect 7728 4664 7866 4990
rect 8392 4800 10064 4838
rect 8392 4790 9984 4800
rect 8392 4738 8450 4790
rect 8502 4748 9984 4790
rect 10036 4748 10064 4800
rect 8502 4738 10064 4748
rect 8392 4698 10064 4738
rect 7728 4612 7767 4664
rect 7819 4612 7866 4664
rect 7728 4600 7866 4612
rect 7728 4548 7767 4600
rect 7819 4548 7866 4600
rect 145 3568 257 3582
rect 145 3482 158 3568
rect 244 3482 257 3568
rect 145 3469 257 3482
rect 5626 3422 6166 3570
rect 232 3209 2153 3326
rect 232 3089 349 3209
rect 64 3079 349 3089
rect 323 2937 349 3079
rect 6062 3158 6166 3422
rect 7728 3242 7866 4548
rect 7364 3158 7490 3160
rect 6062 3127 7490 3158
rect 6062 3071 7397 3127
rect 7453 3071 7490 3127
rect 6062 3048 7490 3071
rect 7364 3046 7490 3048
rect 64 2927 349 2937
rect 7570 3014 7674 3052
rect 7570 2958 7600 3014
rect 7656 2958 7674 3014
rect 6054 2923 6475 2933
rect 7570 2928 7674 2958
rect 6475 2888 7514 2922
rect 6475 2836 7439 2888
rect 7491 2836 7514 2888
rect 6475 2806 7514 2836
rect 6054 2796 6475 2806
rect 7386 2726 7484 2736
rect 7386 2724 7414 2726
rect 7386 2668 7409 2724
rect 7466 2674 7484 2726
rect 7465 2668 7484 2674
rect 7386 2656 7484 2668
rect 7720 2690 7866 3242
rect 8582 3048 8692 3054
rect 8208 3022 8696 3048
rect 8208 3020 8254 3022
rect 8208 2964 8248 3020
rect 8306 3015 8696 3022
rect 8306 2970 8614 3015
rect 8304 2964 8614 2970
rect 8208 2963 8614 2964
rect 8666 2963 8696 3015
rect 8208 2938 8696 2963
rect 9720 2712 9894 2722
rect 7720 2566 9720 2690
rect 7826 2564 9720 2566
rect 147 2539 259 2552
rect 147 2453 159 2539
rect 245 2453 259 2539
rect 147 2439 259 2453
rect 9720 2346 9894 2356
rect 12004 2701 12128 2742
rect 12004 2649 12043 2701
rect 12095 2649 12128 2701
rect 8066 2134 8220 2188
rect 8066 2082 8114 2134
rect 8166 2082 8220 2134
rect 8066 1650 8220 2082
rect 12004 2128 12128 2649
rect 13098 2128 13594 2130
rect 12004 2113 13594 2128
rect 12004 2061 13508 2113
rect 13560 2061 13594 2113
rect 12004 2024 13594 2061
rect 9462 1871 9628 1906
rect 9462 1819 9525 1871
rect 9577 1819 9628 1871
rect 8066 1640 8516 1650
rect 8066 1454 8070 1640
rect 8066 1444 8516 1454
rect 8066 0 8220 1444
rect 9462 1280 9628 1819
rect 9462 1239 11622 1280
rect 9462 1187 11499 1239
rect 11551 1187 11622 1239
rect 9462 1132 11622 1187
<< via2 >>
rect 158 3482 244 3568
rect 7397 3071 7453 3127
rect 7600 3011 7656 3014
rect 7600 2959 7652 3011
rect 7652 2959 7656 3011
rect 7600 2958 7656 2959
rect 6054 2806 6475 2923
rect 7409 2674 7414 2724
rect 7414 2674 7465 2724
rect 7409 2668 7465 2674
rect 8248 2970 8254 3020
rect 8254 2970 8304 3020
rect 8248 2964 8304 2970
rect 159 2453 245 2539
<< metal3 >>
rect 0 5397 2272 5544
rect 145 3573 257 3582
rect 145 3477 153 3573
rect 249 3477 257 3573
rect 145 3469 257 3477
rect 3586 3403 3596 3537
rect 4019 3403 4029 3537
rect 3900 3258 4019 3403
rect 3900 3139 4637 3258
rect 4518 2925 4637 3139
rect 7370 3127 7492 3158
rect 7370 3071 7397 3127
rect 7453 3071 7492 3127
rect 6044 2925 6485 2928
rect 4518 2923 6485 2925
rect 4518 2806 6054 2923
rect 6475 2806 6485 2923
rect 6044 2801 6485 2806
rect 7370 2724 7492 3071
rect 7604 3054 8396 3056
rect 7568 3020 8396 3054
rect 7568 3014 8248 3020
rect 7568 2958 7600 3014
rect 7656 2964 8248 3014
rect 8304 2964 8396 3020
rect 7656 2958 8396 2964
rect 7568 2940 8396 2958
rect 7568 2926 7690 2940
rect 7370 2668 7409 2724
rect 7465 2668 7492 2724
rect 7370 2644 7492 2668
rect 147 2544 259 2552
rect 147 2448 154 2544
rect 250 2448 259 2544
rect 147 2439 259 2448
<< via3 >>
rect 153 3568 249 3573
rect 153 3482 158 3568
rect 158 3482 244 3568
rect 244 3482 249 3568
rect 153 3477 249 3482
rect 3596 3403 4019 3537
rect 154 2539 250 2544
rect 154 2453 159 2539
rect 159 2453 245 2539
rect 245 2453 250 2539
rect 154 2448 250 2453
<< metal4 >>
rect 0 3618 338 3828
rect 152 3573 250 3618
rect 152 3477 153 3573
rect 249 3477 250 3573
rect 3595 3537 4020 3538
rect 3595 3536 3596 3537
rect 152 3476 250 3477
rect 2446 3403 3596 3536
rect 4019 3403 4020 3537
rect 2446 3402 4020 3403
rect 153 2544 251 2545
rect 153 2448 154 2544
rect 250 2448 251 2544
rect 153 2404 251 2448
rect 0 2194 400 2404
use LVDS1  LVDS1_0
timestamp 1699818132
transform 1 0 6383 0 1 3368
box -17 -1584 3470 2114
use LVDS2  LVDS2_0
timestamp 1699818132
transform 1 0 10282 0 1 2832
box -152 -1748 5398 2676
use LVDSBias  LVDSBias_0
timestamp 1699818132
transform 1 0 3502 0 1 5212
box -3498 -5188 2356 652
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0
timestamp 1699818132
transform 1 0 203 0 1 2745
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_1
timestamp 1699818132
transform 1 0 203 0 1 3276
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_2
timestamp 1699818132
transform 1 0 8994 0 1 1512
box -198 -198 198 198
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699818132
transform 1 0 16070 0 1 2446
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1699818132
transform 1 0 16968 0 1 2464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1699818132
transform 1 0 17858 0 1 2480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1699818132
transform 1 0 18884 0 1 2498
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699818132
transform 1 0 19236 0 1 2496
box -38 -48 130 592
<< labels >>
rlabel metal1 s 19252 2582 19290 2624 4 OUT
port 1 nsew
flabel metal3 0 5397 396 5544 0 FreeSans 480 0 0 0 C1
port 2 nsew
flabel metal4 0 3618 338 3828 0 FreeSans 480 0 0 0 INP
port 3 nsew
flabel metal4 0 2194 338 2404 0 FreeSans 480 0 0 0 INN
port 4 nsew
flabel metal2 8066 0 8220 928 0 FreeSans 480 90 0 0 VBIASN
port 5 nsew
flabel metal1 9412 4 19328 1171 0 FreeSans 1600 0 0 0 GND
port 6 nsew
flabel metal1 3372 5570 19328 5860 0 FreeSans 1600 0 0 0 VDD
port 7 nsew
flabel metal1 s 19164 2574 19328 2646 0 FreeSans 480 0 0 0 OUT
port 8 nsew
<< end >>
