magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< pwell >>
rect -175 182 175 216
rect -175 -182 -141 182
rect 141 -182 175 182
rect -175 -216 175 -182
<< nmoslvt >>
rect -15 -42 15 42
<< ndiff >>
rect -73 17 -15 42
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -42 -15 -17
rect 15 17 73 42
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -42 73 -17
<< ndiffc >>
rect -61 -17 -27 17
rect 27 -17 61 17
<< psubdiff >>
rect -175 182 -51 216
rect -17 182 17 216
rect 51 182 175 216
rect -175 119 -141 182
rect -175 51 -141 85
rect 141 119 175 182
rect 141 51 175 85
rect -175 -17 -141 17
rect 141 -17 175 17
rect -175 -85 -141 -51
rect -175 -182 -141 -119
rect 141 -85 175 -51
rect 141 -182 175 -119
rect -175 -216 -51 -182
rect -17 -216 17 -182
rect 51 -216 175 -182
<< psubdiffcont >>
rect -51 182 -17 216
rect 17 182 51 216
rect -175 85 -141 119
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect 141 -119 175 -85
rect -51 -216 -17 -182
rect 17 -216 51 -182
<< poly >>
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -33 64 33 80
rect -15 42 15 64
rect -15 -64 15 -42
rect -33 -80 33 -64
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
<< polycont >>
rect -17 80 17 114
rect -17 -114 17 -80
<< locali >>
rect -175 182 -51 216
rect -17 182 17 216
rect 51 182 175 216
rect -175 119 -141 182
rect 141 119 175 182
rect -175 51 -141 85
rect -33 80 -17 114
rect 17 80 33 114
rect 141 51 175 85
rect -175 -17 -141 17
rect -61 17 -27 46
rect -61 -46 -27 -17
rect 27 17 61 46
rect 27 -46 61 -17
rect 141 -17 175 17
rect -175 -85 -141 -51
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect 141 -85 175 -51
rect -175 -182 -141 -119
rect 141 -182 175 -119
rect -175 -216 -51 -182
rect -17 -216 17 -182
rect 51 -216 175 -182
<< properties >>
string FIXED_BBOX -158 -199 158 199
<< end >>
