VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LVDStop
  CLASS BLOCK ;
  FOREIGN LVDStop ;
  ORIGIN 0.000 0.000 ;
  SIZE 96.830 BY 29.320 ;
  PIN OUT
    ANTENNADIFFAREA 1.287000 ;
    PORT
      LAYER met1 ;
        RECT 95.730 12.870 96.640 13.230 ;
    END
  END OUT
  PIN C1
    ANTENNAGATEAREA 0.442500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.985 11.360 27.720 ;
    END
  END C1
  PIN INP
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met4 ;
        RECT 0.000 18.090 2.560 19.140 ;
    END
  END INP
  PIN INN
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met4 ;
        RECT 0.000 10.970 2.610 12.020 ;
    END
  END INN
  PIN VBIASN
    ANTENNAGATEAREA 45.200001 ;
    ANTENNADIFFAREA 1.810000 ;
    PORT
      LAYER met2 ;
        RECT 40.330 0.000 41.100 7.270 ;
    END
  END VBIASN
  PIN GND
    ANTENNADIFFAREA 69.391800 ;
    PORT
      LAYER met1 ;
        RECT 46.500 0.020 96.640 5.855 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA 102.742401 ;
    PORT
      LAYER met1 ;
        RECT 16.860 27.850 96.640 29.300 ;
    END
  END VDD
  PIN OUT
    PORT
      LAYER met1 ;
        RECT 95.820 12.870 96.640 13.230 ;
    END
  END OUT
  OBS
      LAYER li1 ;
        RECT 0.205 0.120 96.640 29.145 ;
      LAYER met1 ;
        RECT 0.260 27.570 16.580 29.310 ;
        RECT 0.260 13.510 96.640 27.570 ;
        RECT 0.260 12.590 95.450 13.510 ;
        RECT 0.260 6.135 96.640 12.590 ;
        RECT 0.260 0.020 46.220 6.135 ;
      LAYER met2 ;
        RECT 0.320 7.550 77.790 27.705 ;
        RECT 0.320 5.660 40.050 7.550 ;
        RECT 41.380 5.660 77.790 7.550 ;
      LAYER met3 ;
        RECT 11.760 26.585 41.980 27.755 ;
        RECT 0.725 9.320 41.980 26.585 ;
      LAYER met4 ;
        RECT 0.760 19.540 28.900 23.270 ;
        RECT 2.960 17.690 28.900 19.540 ;
        RECT 0.760 12.420 28.900 17.690 ;
        RECT 3.010 10.570 28.900 12.420 ;
        RECT 0.760 9.380 28.900 10.570 ;
  END
END LVDStop
END LIBRARY

