magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< nwell >>
rect -348 312 118 652
<< psubdiff >>
rect -358 23 -334 94
rect -212 23 -188 94
<< nsubdiff >>
rect -303 501 -161 534
rect -303 413 -274 501
rect -191 413 -161 501
rect -303 387 -161 413
<< psubdiffcont >>
rect -334 23 -212 94
<< nsubdiffcont >>
rect -274 413 -191 501
<< locali >>
rect -297 501 -169 527
rect -297 413 -274 501
rect -191 413 -169 501
rect -297 388 -169 413
rect 88 324 92 358
rect 126 324 130 358
rect 226 324 230 358
rect 264 324 268 358
rect 402 324 406 358
rect 440 324 444 358
rect -523 278 -522 312
rect 164 209 340 237
rect 238 128 272 156
rect -387 23 -334 94
rect -212 23 -196 94
rect 512 13 632 354
rect 764 324 768 358
rect 802 324 806 358
rect 878 324 882 358
rect 916 324 920 358
rect 1008 324 1012 358
rect 1046 324 1050 358
rect 801 210 977 235
rect 902 127 938 158
rect -1042 -257 -972 -238
rect -1042 -291 -1024 -257
rect -990 -291 -972 -257
rect -1042 -329 -972 -291
rect -1042 -363 -1024 -329
rect -990 -363 -972 -329
rect -1042 -401 -972 -363
rect -1042 -435 -1024 -401
rect -990 -435 -972 -401
rect -1042 -473 -972 -435
rect -1042 -507 -1024 -473
rect -990 -507 -972 -473
rect -1042 -545 -972 -507
rect -1042 -579 -1024 -545
rect -990 -579 -972 -545
rect -1042 -617 -972 -579
rect -1042 -651 -1024 -617
rect -990 -651 -972 -617
rect -1042 -670 -972 -651
rect -724 -257 -654 -238
rect -724 -291 -706 -257
rect -672 -291 -654 -257
rect -724 -329 -654 -291
rect -724 -363 -706 -329
rect -672 -363 -654 -329
rect -724 -401 -654 -363
rect -724 -435 -706 -401
rect -672 -435 -654 -401
rect -724 -473 -654 -435
rect -724 -507 -706 -473
rect -672 -507 -654 -473
rect -724 -545 -654 -507
rect -724 -579 -706 -545
rect -672 -579 -654 -545
rect -724 -617 -654 -579
rect -724 -651 -706 -617
rect -672 -651 -654 -617
rect -724 -670 -654 -651
rect -406 -257 -336 -238
rect -406 -291 -388 -257
rect -354 -291 -336 -257
rect -406 -329 -336 -291
rect -406 -363 -388 -329
rect -354 -363 -336 -329
rect -406 -401 -336 -363
rect -406 -435 -388 -401
rect -354 -435 -336 -401
rect -406 -473 -336 -435
rect -406 -507 -388 -473
rect -354 -507 -336 -473
rect -406 -545 -336 -507
rect -406 -579 -388 -545
rect -354 -579 -336 -545
rect -406 -617 -336 -579
rect -406 -651 -388 -617
rect -354 -651 -336 -617
rect -406 -670 -336 -651
rect -88 -257 -18 -238
rect -88 -291 -70 -257
rect -36 -291 -18 -257
rect -88 -329 -18 -291
rect -88 -363 -70 -329
rect -36 -363 -18 -329
rect -88 -401 -18 -363
rect -88 -435 -70 -401
rect -36 -435 -18 -401
rect -88 -473 -18 -435
rect -88 -507 -70 -473
rect -36 -507 -18 -473
rect -88 -545 -18 -507
rect -88 -579 -70 -545
rect -36 -579 -18 -545
rect -88 -617 -18 -579
rect -88 -651 -70 -617
rect -36 -651 -18 -617
rect -88 -670 -18 -651
rect 230 -257 300 -238
rect 230 -291 248 -257
rect 282 -291 300 -257
rect 230 -329 300 -291
rect 230 -363 248 -329
rect 282 -363 300 -329
rect 230 -401 300 -363
rect 230 -435 248 -401
rect 282 -435 300 -401
rect 230 -473 300 -435
rect 230 -507 248 -473
rect 282 -507 300 -473
rect 230 -545 300 -507
rect 230 -579 248 -545
rect 282 -579 300 -545
rect 230 -617 300 -579
rect 230 -651 248 -617
rect 282 -651 300 -617
rect 230 -670 300 -651
rect -1042 -1089 -972 -1070
rect -1042 -1123 -1024 -1089
rect -990 -1123 -972 -1089
rect -1042 -1161 -972 -1123
rect -1042 -1195 -1024 -1161
rect -990 -1195 -972 -1161
rect -1042 -1233 -972 -1195
rect -1042 -1267 -1024 -1233
rect -990 -1267 -972 -1233
rect -1042 -1305 -972 -1267
rect -1042 -1339 -1024 -1305
rect -990 -1339 -972 -1305
rect -1042 -1377 -972 -1339
rect -1042 -1411 -1024 -1377
rect -990 -1411 -972 -1377
rect -1042 -1449 -972 -1411
rect -1042 -1483 -1024 -1449
rect -990 -1483 -972 -1449
rect -1042 -1502 -972 -1483
rect -724 -1089 -654 -1070
rect -724 -1123 -706 -1089
rect -672 -1123 -654 -1089
rect -724 -1161 -654 -1123
rect -724 -1195 -706 -1161
rect -672 -1195 -654 -1161
rect -724 -1233 -654 -1195
rect -724 -1267 -706 -1233
rect -672 -1267 -654 -1233
rect -724 -1305 -654 -1267
rect -724 -1339 -706 -1305
rect -672 -1339 -654 -1305
rect -724 -1377 -654 -1339
rect -724 -1411 -706 -1377
rect -672 -1411 -654 -1377
rect -724 -1449 -654 -1411
rect -724 -1483 -706 -1449
rect -672 -1483 -654 -1449
rect -724 -1502 -654 -1483
rect -406 -1089 -336 -1070
rect -406 -1123 -388 -1089
rect -354 -1123 -336 -1089
rect -406 -1161 -336 -1123
rect -406 -1195 -388 -1161
rect -354 -1195 -336 -1161
rect -406 -1233 -336 -1195
rect -406 -1267 -388 -1233
rect -354 -1267 -336 -1233
rect -406 -1305 -336 -1267
rect -406 -1339 -388 -1305
rect -354 -1339 -336 -1305
rect -406 -1377 -336 -1339
rect -406 -1411 -388 -1377
rect -354 -1411 -336 -1377
rect -406 -1449 -336 -1411
rect -406 -1483 -388 -1449
rect -354 -1483 -336 -1449
rect -406 -1502 -336 -1483
rect -88 -1089 -18 -1070
rect -88 -1123 -70 -1089
rect -36 -1123 -18 -1089
rect -88 -1161 -18 -1123
rect -88 -1195 -70 -1161
rect -36 -1195 -18 -1161
rect -88 -1233 -18 -1195
rect -88 -1267 -70 -1233
rect -36 -1267 -18 -1233
rect -88 -1305 -18 -1267
rect -88 -1339 -70 -1305
rect -36 -1339 -18 -1305
rect -88 -1377 -18 -1339
rect -88 -1411 -70 -1377
rect -36 -1411 -18 -1377
rect -88 -1449 -18 -1411
rect -88 -1483 -70 -1449
rect -36 -1483 -18 -1449
rect -88 -1502 -18 -1483
rect 230 -1089 300 -1070
rect 230 -1123 248 -1089
rect 282 -1123 300 -1089
rect 230 -1161 300 -1123
rect 230 -1195 248 -1161
rect 282 -1195 300 -1161
rect 230 -1233 300 -1195
rect 230 -1267 248 -1233
rect 282 -1267 300 -1233
rect 230 -1305 300 -1267
rect 230 -1339 248 -1305
rect 282 -1339 300 -1305
rect 230 -1377 300 -1339
rect 230 -1411 248 -1377
rect 282 -1411 300 -1377
rect 230 -1449 300 -1411
rect 230 -1483 248 -1449
rect 282 -1483 300 -1449
rect 230 -1502 300 -1483
rect -720 -1600 -662 -1596
rect -720 -1609 -708 -1600
rect -1154 -1634 -708 -1609
rect -674 -1609 -662 -1600
rect -674 -1634 -510 -1609
rect 405 -1624 770 -104
rect 884 -253 954 -234
rect 884 -287 902 -253
rect 936 -287 954 -253
rect 884 -325 954 -287
rect 884 -359 902 -325
rect 936 -359 954 -325
rect 884 -397 954 -359
rect 884 -431 902 -397
rect 936 -431 954 -397
rect 884 -469 954 -431
rect 884 -503 902 -469
rect 936 -503 954 -469
rect 884 -541 954 -503
rect 884 -575 902 -541
rect 936 -575 954 -541
rect 884 -613 954 -575
rect 884 -647 902 -613
rect 936 -647 954 -613
rect 884 -666 954 -647
rect 1202 -253 1272 -234
rect 1202 -287 1220 -253
rect 1254 -287 1272 -253
rect 1202 -325 1272 -287
rect 1202 -359 1220 -325
rect 1254 -359 1272 -325
rect 1202 -397 1272 -359
rect 1202 -431 1220 -397
rect 1254 -431 1272 -397
rect 1202 -469 1272 -431
rect 1202 -503 1220 -469
rect 1254 -503 1272 -469
rect 1202 -541 1272 -503
rect 1202 -575 1220 -541
rect 1254 -575 1272 -541
rect 1202 -613 1272 -575
rect 1202 -647 1220 -613
rect 1254 -647 1272 -613
rect 1202 -666 1272 -647
rect 1520 -253 1590 -234
rect 1520 -287 1538 -253
rect 1572 -287 1590 -253
rect 1520 -325 1590 -287
rect 1520 -359 1538 -325
rect 1572 -359 1590 -325
rect 1520 -397 1590 -359
rect 1520 -431 1538 -397
rect 1572 -431 1590 -397
rect 1520 -469 1590 -431
rect 1520 -503 1538 -469
rect 1572 -503 1590 -469
rect 1520 -541 1590 -503
rect 1520 -575 1538 -541
rect 1572 -575 1590 -541
rect 1520 -613 1590 -575
rect 1520 -647 1538 -613
rect 1572 -647 1590 -613
rect 1520 -666 1590 -647
rect 1838 -253 1908 -234
rect 1838 -287 1856 -253
rect 1890 -287 1908 -253
rect 1838 -325 1908 -287
rect 1838 -359 1856 -325
rect 1890 -359 1908 -325
rect 1838 -397 1908 -359
rect 1838 -431 1856 -397
rect 1890 -431 1908 -397
rect 1838 -469 1908 -431
rect 1838 -503 1856 -469
rect 1890 -503 1908 -469
rect 1838 -541 1908 -503
rect 1838 -575 1856 -541
rect 1890 -575 1908 -541
rect 1838 -613 1908 -575
rect 1838 -647 1856 -613
rect 1890 -647 1908 -613
rect 1838 -666 1908 -647
rect 2156 -253 2226 -234
rect 2156 -287 2174 -253
rect 2208 -287 2226 -253
rect 2156 -325 2226 -287
rect 2156 -359 2174 -325
rect 2208 -359 2226 -325
rect 2156 -397 2226 -359
rect 2156 -431 2174 -397
rect 2208 -431 2226 -397
rect 2156 -469 2226 -431
rect 2156 -503 2174 -469
rect 2208 -503 2226 -469
rect 2156 -541 2226 -503
rect 2156 -575 2174 -541
rect 2208 -575 2226 -541
rect 2156 -613 2226 -575
rect 2156 -647 2174 -613
rect 2208 -647 2226 -613
rect 2156 -666 2226 -647
rect 884 -1085 954 -1066
rect 884 -1119 902 -1085
rect 936 -1119 954 -1085
rect 884 -1157 954 -1119
rect 884 -1191 902 -1157
rect 936 -1191 954 -1157
rect 884 -1229 954 -1191
rect 884 -1263 902 -1229
rect 936 -1263 954 -1229
rect 884 -1301 954 -1263
rect 884 -1335 902 -1301
rect 936 -1335 954 -1301
rect 884 -1373 954 -1335
rect 884 -1407 902 -1373
rect 936 -1407 954 -1373
rect 884 -1445 954 -1407
rect 884 -1479 902 -1445
rect 936 -1479 954 -1445
rect 884 -1498 954 -1479
rect 1202 -1085 1272 -1066
rect 1202 -1119 1220 -1085
rect 1254 -1119 1272 -1085
rect 1202 -1157 1272 -1119
rect 1202 -1191 1220 -1157
rect 1254 -1191 1272 -1157
rect 1202 -1229 1272 -1191
rect 1202 -1263 1220 -1229
rect 1254 -1263 1272 -1229
rect 1202 -1301 1272 -1263
rect 1202 -1335 1220 -1301
rect 1254 -1335 1272 -1301
rect 1202 -1373 1272 -1335
rect 1202 -1407 1220 -1373
rect 1254 -1407 1272 -1373
rect 1202 -1445 1272 -1407
rect 1202 -1479 1220 -1445
rect 1254 -1479 1272 -1445
rect 1202 -1498 1272 -1479
rect 1520 -1085 1590 -1066
rect 1520 -1119 1538 -1085
rect 1572 -1119 1590 -1085
rect 1520 -1157 1590 -1119
rect 1520 -1191 1538 -1157
rect 1572 -1191 1590 -1157
rect 1520 -1229 1590 -1191
rect 1520 -1263 1538 -1229
rect 1572 -1263 1590 -1229
rect 1520 -1301 1590 -1263
rect 1520 -1335 1538 -1301
rect 1572 -1335 1590 -1301
rect 1520 -1373 1590 -1335
rect 1520 -1407 1538 -1373
rect 1572 -1407 1590 -1373
rect 1520 -1445 1590 -1407
rect 1520 -1479 1538 -1445
rect 1572 -1479 1590 -1445
rect 1520 -1498 1590 -1479
rect 1838 -1085 1908 -1066
rect 1838 -1119 1856 -1085
rect 1890 -1119 1908 -1085
rect 1838 -1157 1908 -1119
rect 1838 -1191 1856 -1157
rect 1890 -1191 1908 -1157
rect 1838 -1229 1908 -1191
rect 1838 -1263 1856 -1229
rect 1890 -1263 1908 -1229
rect 1838 -1301 1908 -1263
rect 1838 -1335 1856 -1301
rect 1890 -1335 1908 -1301
rect 1838 -1373 1908 -1335
rect 1838 -1407 1856 -1373
rect 1890 -1407 1908 -1373
rect 1838 -1445 1908 -1407
rect 1838 -1479 1856 -1445
rect 1890 -1479 1908 -1445
rect 1838 -1498 1908 -1479
rect 2156 -1085 2226 -1066
rect 2156 -1119 2174 -1085
rect 2208 -1119 2226 -1085
rect 2156 -1157 2226 -1119
rect 2156 -1191 2174 -1157
rect 2208 -1191 2226 -1157
rect 2156 -1229 2226 -1191
rect 2156 -1263 2174 -1229
rect 2208 -1263 2226 -1229
rect 2156 -1301 2226 -1263
rect 2156 -1335 2174 -1301
rect 2208 -1335 2226 -1301
rect 2156 -1373 2226 -1335
rect 2156 -1407 2174 -1373
rect 2208 -1407 2226 -1373
rect 2156 -1445 2226 -1407
rect 2156 -1479 2174 -1445
rect 2208 -1479 2226 -1445
rect 2156 -1498 2226 -1479
rect 1838 -1592 1896 -1588
rect 1838 -1601 1850 -1592
rect -1154 -1862 -510 -1634
rect 1720 -1626 1850 -1601
rect 1884 -1601 1896 -1592
rect 1884 -1626 2354 -1601
rect 1720 -1810 2354 -1626
rect 1720 -1837 1848 -1810
rect 1836 -1844 1848 -1837
rect 1882 -1837 2354 -1810
rect 1882 -1844 1894 -1837
rect 1836 -1848 1894 -1844
rect -1154 -1872 -712 -1862
rect -724 -1896 -712 -1872
rect -678 -1872 -510 -1862
rect -678 -1896 -666 -1872
rect -724 -1900 -666 -1896
rect 1834 -1959 1904 -1940
rect 1834 -1993 1852 -1959
rect 1886 -1993 1904 -1959
rect -1030 -2013 -960 -1994
rect -1030 -2047 -1012 -2013
rect -978 -2047 -960 -2013
rect -1030 -2085 -960 -2047
rect -1030 -2119 -1012 -2085
rect -978 -2119 -960 -2085
rect -1030 -2157 -960 -2119
rect -1030 -2191 -1012 -2157
rect -978 -2191 -960 -2157
rect -1030 -2229 -960 -2191
rect -1030 -2263 -1012 -2229
rect -978 -2263 -960 -2229
rect -1030 -2301 -960 -2263
rect -1030 -2335 -1012 -2301
rect -978 -2335 -960 -2301
rect -1030 -2373 -960 -2335
rect -1030 -2407 -1012 -2373
rect -978 -2407 -960 -2373
rect -1030 -2426 -960 -2407
rect -712 -2013 -642 -1994
rect -712 -2047 -694 -2013
rect -660 -2047 -642 -2013
rect -712 -2085 -642 -2047
rect -712 -2119 -694 -2085
rect -660 -2119 -642 -2085
rect -712 -2157 -642 -2119
rect -712 -2191 -694 -2157
rect -660 -2191 -642 -2157
rect -712 -2229 -642 -2191
rect -712 -2263 -694 -2229
rect -660 -2263 -642 -2229
rect -712 -2301 -642 -2263
rect -712 -2335 -694 -2301
rect -660 -2335 -642 -2301
rect -712 -2373 -642 -2335
rect 1834 -2031 1904 -1993
rect 1834 -2065 1852 -2031
rect 1886 -2065 1904 -2031
rect 1834 -2103 1904 -2065
rect 1834 -2137 1852 -2103
rect 1886 -2137 1904 -2103
rect 1834 -2175 1904 -2137
rect 1834 -2209 1852 -2175
rect 1886 -2209 1904 -2175
rect 1834 -2247 1904 -2209
rect 1834 -2281 1852 -2247
rect 1886 -2281 1904 -2247
rect 1834 -2319 1904 -2281
rect 1834 -2353 1852 -2319
rect 1886 -2353 1904 -2319
rect 1834 -2372 1904 -2353
rect 2152 -1959 2222 -1940
rect 2152 -1993 2170 -1959
rect 2204 -1993 2222 -1959
rect 2152 -2031 2222 -1993
rect 2152 -2065 2170 -2031
rect 2204 -2065 2222 -2031
rect 2152 -2103 2222 -2065
rect 2152 -2137 2170 -2103
rect 2204 -2137 2222 -2103
rect 2152 -2175 2222 -2137
rect 2152 -2209 2170 -2175
rect 2204 -2209 2222 -2175
rect 2152 -2247 2222 -2209
rect 2152 -2281 2170 -2247
rect 2204 -2281 2222 -2247
rect 2152 -2319 2222 -2281
rect 2152 -2353 2170 -2319
rect 2204 -2353 2222 -2319
rect 2152 -2372 2222 -2353
rect -712 -2407 -694 -2373
rect -660 -2407 -642 -2373
rect -712 -2426 -642 -2407
rect -523 -2770 -403 -2493
rect 1370 -2596 1408 -2562
rect -198 -2638 -160 -2604
rect 1370 -2684 1408 -2650
rect -198 -2726 -160 -2692
rect -548 -2771 -403 -2770
rect -548 -2805 -547 -2771
rect -513 -2805 -403 -2771
rect 1246 -2765 1304 -2764
rect 1246 -2799 1258 -2765
rect 1292 -2799 1304 -2765
rect 1246 -2800 1304 -2799
rect 1370 -2765 1428 -2764
rect 1370 -2799 1382 -2765
rect 1416 -2799 1428 -2765
rect 1370 -2800 1428 -2799
rect 1474 -2765 1532 -2764
rect 1474 -2799 1486 -2765
rect 1520 -2799 1532 -2765
rect 1606 -2788 1726 -2450
rect 1606 -2789 1738 -2788
rect 1606 -2791 1703 -2789
rect 1474 -2800 1532 -2799
rect -548 -2806 -403 -2805
rect -523 -2812 -403 -2806
rect -544 -2860 -403 -2812
rect -322 -2805 -264 -2804
rect -322 -2839 -310 -2805
rect -276 -2839 -264 -2805
rect -94 -2805 -36 -2804
rect -322 -2840 -264 -2839
rect -206 -2807 -148 -2806
rect -206 -2841 -194 -2807
rect -160 -2841 -148 -2807
rect -94 -2839 -82 -2805
rect -48 -2839 -36 -2805
rect 1702 -2823 1703 -2791
rect 1737 -2823 1738 -2789
rect 1702 -2824 1738 -2823
rect -94 -2840 -36 -2839
rect -206 -2842 -148 -2841
rect -546 -2861 -403 -2860
rect -546 -2895 -545 -2861
rect -511 -2895 -403 -2861
rect -546 -2896 -403 -2895
rect -544 -2901 -403 -2896
rect 1702 -2863 1738 -2862
rect 1702 -2897 1703 -2863
rect 1737 -2897 1738 -2863
rect 1702 -2898 1738 -2897
rect 1834 -4591 1904 -4572
rect 1834 -4625 1852 -4591
rect 1886 -4625 1904 -4591
rect -1030 -4645 -960 -4626
rect -1030 -4679 -1012 -4645
rect -978 -4679 -960 -4645
rect -1030 -4717 -960 -4679
rect -1030 -4751 -1012 -4717
rect -978 -4751 -960 -4717
rect -1030 -4789 -960 -4751
rect -1030 -4823 -1012 -4789
rect -978 -4823 -960 -4789
rect -1030 -4861 -960 -4823
rect -1030 -4895 -1012 -4861
rect -978 -4895 -960 -4861
rect -1030 -4933 -960 -4895
rect -1030 -4967 -1012 -4933
rect -978 -4967 -960 -4933
rect -1030 -5005 -960 -4967
rect -1030 -5039 -1012 -5005
rect -978 -5039 -960 -5005
rect -1030 -5058 -960 -5039
rect -712 -4645 -642 -4626
rect -712 -4679 -694 -4645
rect -660 -4679 -642 -4645
rect -712 -4717 -642 -4679
rect -712 -4751 -694 -4717
rect -660 -4751 -642 -4717
rect -712 -4789 -642 -4751
rect -712 -4823 -694 -4789
rect -660 -4823 -642 -4789
rect -712 -4861 -642 -4823
rect -712 -4895 -694 -4861
rect -660 -4895 -642 -4861
rect -712 -4933 -642 -4895
rect -712 -4967 -694 -4933
rect -660 -4967 -642 -4933
rect -712 -5005 -642 -4967
rect 1834 -4663 1904 -4625
rect 1834 -4697 1852 -4663
rect 1886 -4697 1904 -4663
rect 1834 -4735 1904 -4697
rect 1834 -4769 1852 -4735
rect 1886 -4769 1904 -4735
rect 1834 -4807 1904 -4769
rect 1834 -4841 1852 -4807
rect 1886 -4841 1904 -4807
rect 1834 -4879 1904 -4841
rect 1834 -4913 1852 -4879
rect 1886 -4913 1904 -4879
rect 1834 -4951 1904 -4913
rect 1834 -4985 1852 -4951
rect 1886 -4985 1904 -4951
rect 1834 -5004 1904 -4985
rect 2152 -4591 2222 -4572
rect 2152 -4625 2170 -4591
rect 2204 -4625 2222 -4591
rect 2152 -4663 2222 -4625
rect 2152 -4697 2170 -4663
rect 2204 -4697 2222 -4663
rect 2152 -4735 2222 -4697
rect 2152 -4769 2170 -4735
rect 2204 -4769 2222 -4735
rect 2152 -4807 2222 -4769
rect 2152 -4841 2170 -4807
rect 2204 -4841 2222 -4807
rect 2152 -4879 2222 -4841
rect 2152 -4913 2170 -4879
rect 2204 -4913 2222 -4879
rect 2152 -4951 2222 -4913
rect 2152 -4985 2170 -4951
rect 2204 -4985 2222 -4951
rect 2152 -5004 2222 -4985
rect -712 -5039 -694 -5005
rect -660 -5039 -642 -5005
rect -712 -5058 -642 -5039
<< viali >>
rect -274 413 -191 501
rect 92 324 126 358
rect 230 324 264 358
rect 406 324 440 358
rect -659 271 -523 319
rect -460 213 -324 261
rect 156 237 348 279
rect 71 165 105 199
rect 399 165 433 199
rect -334 23 -212 94
rect 156 86 348 128
rect 768 324 802 358
rect 882 324 916 358
rect 1012 324 1046 358
rect 795 235 987 277
rect 708 166 742 200
rect 1051 149 1088 216
rect 792 85 984 127
rect -1024 -291 -990 -257
rect -1024 -363 -990 -329
rect -1024 -435 -990 -401
rect -1024 -507 -990 -473
rect -1024 -579 -990 -545
rect -1024 -651 -990 -617
rect -706 -291 -672 -257
rect -706 -363 -672 -329
rect -706 -435 -672 -401
rect -706 -507 -672 -473
rect -706 -579 -672 -545
rect -706 -651 -672 -617
rect -388 -291 -354 -257
rect -388 -363 -354 -329
rect -388 -435 -354 -401
rect -388 -507 -354 -473
rect -388 -579 -354 -545
rect -388 -651 -354 -617
rect -70 -291 -36 -257
rect -70 -363 -36 -329
rect -70 -435 -36 -401
rect -70 -507 -36 -473
rect -70 -579 -36 -545
rect -70 -651 -36 -617
rect 248 -291 282 -257
rect 248 -363 282 -329
rect 248 -435 282 -401
rect 248 -507 282 -473
rect 248 -579 282 -545
rect 248 -651 282 -617
rect -1024 -1123 -990 -1089
rect -1024 -1195 -990 -1161
rect -1024 -1267 -990 -1233
rect -1024 -1339 -990 -1305
rect -1024 -1411 -990 -1377
rect -1024 -1483 -990 -1449
rect -706 -1123 -672 -1089
rect -706 -1195 -672 -1161
rect -706 -1267 -672 -1233
rect -706 -1339 -672 -1305
rect -706 -1411 -672 -1377
rect -706 -1483 -672 -1449
rect -388 -1123 -354 -1089
rect -388 -1195 -354 -1161
rect -388 -1267 -354 -1233
rect -388 -1339 -354 -1305
rect -388 -1411 -354 -1377
rect -388 -1483 -354 -1449
rect -70 -1123 -36 -1089
rect -70 -1195 -36 -1161
rect -70 -1267 -36 -1233
rect -70 -1339 -36 -1305
rect -70 -1411 -36 -1377
rect -70 -1483 -36 -1449
rect 248 -1123 282 -1089
rect 248 -1195 282 -1161
rect 248 -1267 282 -1233
rect 248 -1339 282 -1305
rect 248 -1411 282 -1377
rect 248 -1483 282 -1449
rect -708 -1634 -674 -1600
rect 902 -287 936 -253
rect 902 -359 936 -325
rect 902 -431 936 -397
rect 902 -503 936 -469
rect 902 -575 936 -541
rect 902 -647 936 -613
rect 1220 -287 1254 -253
rect 1220 -359 1254 -325
rect 1220 -431 1254 -397
rect 1220 -503 1254 -469
rect 1220 -575 1254 -541
rect 1220 -647 1254 -613
rect 1538 -287 1572 -253
rect 1538 -359 1572 -325
rect 1538 -431 1572 -397
rect 1538 -503 1572 -469
rect 1538 -575 1572 -541
rect 1538 -647 1572 -613
rect 1856 -287 1890 -253
rect 1856 -359 1890 -325
rect 1856 -431 1890 -397
rect 1856 -503 1890 -469
rect 1856 -575 1890 -541
rect 1856 -647 1890 -613
rect 2174 -287 2208 -253
rect 2174 -359 2208 -325
rect 2174 -431 2208 -397
rect 2174 -503 2208 -469
rect 2174 -575 2208 -541
rect 2174 -647 2208 -613
rect 902 -1119 936 -1085
rect 902 -1191 936 -1157
rect 902 -1263 936 -1229
rect 902 -1335 936 -1301
rect 902 -1407 936 -1373
rect 902 -1479 936 -1445
rect 1220 -1119 1254 -1085
rect 1220 -1191 1254 -1157
rect 1220 -1263 1254 -1229
rect 1220 -1335 1254 -1301
rect 1220 -1407 1254 -1373
rect 1220 -1479 1254 -1445
rect 1538 -1119 1572 -1085
rect 1538 -1191 1572 -1157
rect 1538 -1263 1572 -1229
rect 1538 -1335 1572 -1301
rect 1538 -1407 1572 -1373
rect 1538 -1479 1572 -1445
rect 1856 -1119 1890 -1085
rect 1856 -1191 1890 -1157
rect 1856 -1263 1890 -1229
rect 1856 -1335 1890 -1301
rect 1856 -1407 1890 -1373
rect 1856 -1479 1890 -1445
rect 2174 -1119 2208 -1085
rect 2174 -1191 2208 -1157
rect 2174 -1263 2208 -1229
rect 2174 -1335 2208 -1301
rect 2174 -1407 2208 -1373
rect 2174 -1479 2208 -1445
rect 1850 -1626 1884 -1592
rect 1848 -1844 1882 -1810
rect -712 -1896 -678 -1862
rect 1852 -1993 1886 -1959
rect -1012 -2047 -978 -2013
rect -1012 -2119 -978 -2085
rect -1012 -2191 -978 -2157
rect -1012 -2263 -978 -2229
rect -1012 -2335 -978 -2301
rect -1012 -2407 -978 -2373
rect -694 -2047 -660 -2013
rect -694 -2119 -660 -2085
rect -694 -2191 -660 -2157
rect -694 -2263 -660 -2229
rect -694 -2335 -660 -2301
rect 1852 -2065 1886 -2031
rect 1852 -2137 1886 -2103
rect 1852 -2209 1886 -2175
rect 1852 -2281 1886 -2247
rect 1852 -2353 1886 -2319
rect 2170 -1993 2204 -1959
rect 2170 -2065 2204 -2031
rect 2170 -2137 2204 -2103
rect 2170 -2209 2204 -2175
rect 2170 -2281 2204 -2247
rect 2170 -2353 2204 -2319
rect -694 -2407 -660 -2373
rect 1336 -2596 1370 -2562
rect 1408 -2596 1442 -2562
rect -232 -2638 -198 -2604
rect -160 -2638 -126 -2604
rect 1248 -2640 1282 -2606
rect -72 -2682 -38 -2648
rect 1336 -2684 1370 -2650
rect 1408 -2684 1442 -2650
rect -232 -2726 -198 -2692
rect -160 -2726 -126 -2692
rect -547 -2805 -513 -2771
rect 1258 -2799 1292 -2765
rect 1382 -2799 1416 -2765
rect 1486 -2799 1520 -2765
rect -310 -2839 -276 -2805
rect -194 -2841 -160 -2807
rect -82 -2839 -48 -2805
rect 1703 -2823 1737 -2789
rect -545 -2895 -511 -2861
rect 1703 -2897 1737 -2863
rect 1852 -4625 1886 -4591
rect -1012 -4679 -978 -4645
rect -1012 -4751 -978 -4717
rect -1012 -4823 -978 -4789
rect -1012 -4895 -978 -4861
rect -1012 -4967 -978 -4933
rect -1012 -5039 -978 -5005
rect -694 -4679 -660 -4645
rect -694 -4751 -660 -4717
rect -694 -4823 -660 -4789
rect -694 -4895 -660 -4861
rect -694 -4967 -660 -4933
rect 1852 -4697 1886 -4663
rect 1852 -4769 1886 -4735
rect 1852 -4841 1886 -4807
rect 1852 -4913 1886 -4879
rect 1852 -4985 1886 -4951
rect 2170 -4625 2204 -4591
rect 2170 -4697 2204 -4663
rect 2170 -4769 2204 -4735
rect 2170 -4841 2204 -4807
rect 2170 -4913 2204 -4879
rect 2170 -4985 2204 -4951
rect -694 -5039 -660 -5005
<< metal1 >>
rect -65 648 1228 650
rect -382 552 1228 648
rect -297 501 1228 552
rect -297 413 -274 501
rect -191 413 1228 501
rect -297 388 1228 413
rect -130 358 1228 388
rect -675 320 -502 327
rect -1223 319 -502 320
rect -1234 224 -1224 319
rect -893 271 -659 319
rect -523 271 -502 319
rect -130 324 92 358
rect 126 324 230 358
rect 264 324 406 358
rect 440 324 768 358
rect 802 324 882 358
rect 916 324 1012 358
rect 1046 324 1228 358
rect -130 300 1228 324
rect -893 256 -502 271
rect 144 279 360 300
rect -472 266 -312 268
rect -472 261 -80 266
rect -893 224 -883 256
rect -472 213 -460 261
rect -324 216 -80 261
rect 144 237 156 279
rect 348 237 360 279
rect 144 231 360 237
rect 783 277 999 300
rect 783 235 795 277
rect 987 235 999 277
rect 783 229 999 235
rect 1045 216 1094 228
rect -324 213 112 216
rect -472 206 112 213
rect -130 200 112 206
rect 386 200 749 216
rect 1045 200 1051 216
rect -130 199 708 200
rect -130 165 71 199
rect 105 165 399 199
rect 433 166 708 199
rect 742 166 1051 200
rect 433 165 1051 166
rect -130 164 1051 165
rect -130 142 112 164
rect 386 150 749 164
rect 1045 149 1051 164
rect 1088 149 1094 216
rect 1045 137 1094 149
rect 144 128 360 134
rect -924 90 -631 107
rect -924 21 -903 90
rect -688 21 -631 90
rect -387 94 -186 105
rect -624 83 -572 84
rect -624 30 -572 31
rect -924 9 -631 21
rect -387 23 -334 94
rect -212 23 -186 94
rect 144 86 156 128
rect 348 86 360 128
rect 144 80 360 86
rect 780 127 996 133
rect 780 85 792 127
rect 984 85 996 127
rect -387 8 -186 23
rect -1070 -257 -624 -220
rect -1070 -291 -1024 -257
rect -990 -291 -706 -257
rect -672 -291 -624 -257
rect -1070 -329 -624 -291
rect -1070 -363 -1024 -329
rect -990 -363 -706 -329
rect -672 -363 -624 -329
rect -1070 -401 -624 -363
rect -1070 -435 -1024 -401
rect -990 -435 -706 -401
rect -672 -435 -624 -401
rect -1070 -473 -624 -435
rect -1070 -507 -1024 -473
rect -990 -507 -706 -473
rect -672 -507 -624 -473
rect -1070 -545 -624 -507
rect -1070 -579 -1024 -545
rect -990 -579 -706 -545
rect -672 -579 -624 -545
rect -1070 -617 -624 -579
rect -1070 -651 -1024 -617
rect -990 -651 -706 -617
rect -672 -651 -624 -617
rect -1070 -682 -624 -651
rect -442 -257 8 -206
rect -442 -291 -388 -257
rect -354 -291 -70 -257
rect -36 -291 8 -257
rect -442 -329 8 -291
rect -442 -363 -388 -329
rect -354 -363 -70 -329
rect -36 -363 8 -329
rect -442 -401 8 -363
rect -442 -435 -388 -401
rect -354 -435 -70 -401
rect -36 -435 8 -401
rect -442 -473 8 -435
rect -442 -507 -388 -473
rect -354 -507 -70 -473
rect -36 -507 8 -473
rect -442 -545 8 -507
rect -442 -579 -388 -545
rect -354 -579 -70 -545
rect -36 -579 8 -545
rect -442 -617 8 -579
rect -442 -651 -388 -617
rect -354 -651 -70 -617
rect -36 -651 8 -617
rect -442 -678 8 -651
rect 214 -257 310 80
rect 780 79 996 85
rect 214 -291 248 -257
rect 282 -291 310 -257
rect 214 -329 310 -291
rect 214 -363 248 -329
rect 282 -363 310 -329
rect 214 -401 310 -363
rect 214 -435 248 -401
rect 282 -435 310 -401
rect 214 -473 310 -435
rect 214 -507 248 -473
rect 282 -507 310 -473
rect 214 -545 310 -507
rect 214 -579 248 -545
rect 282 -579 310 -545
rect 214 -617 310 -579
rect 214 -651 248 -617
rect 282 -651 310 -617
rect 214 -684 310 -651
rect 862 -253 968 79
rect 862 -287 902 -253
rect 936 -287 968 -253
rect 862 -325 968 -287
rect 862 -359 902 -325
rect 936 -359 968 -325
rect 862 -397 968 -359
rect 862 -431 902 -397
rect 936 -431 968 -397
rect 862 -469 968 -431
rect 862 -503 902 -469
rect 936 -503 968 -469
rect 862 -541 968 -503
rect 862 -575 902 -541
rect 936 -575 968 -541
rect 862 -613 968 -575
rect 862 -647 902 -613
rect 936 -647 968 -613
rect 862 -676 968 -647
rect 1184 -253 1614 -198
rect 1184 -287 1220 -253
rect 1254 -287 1538 -253
rect 1572 -287 1614 -253
rect 1184 -325 1614 -287
rect 1184 -359 1220 -325
rect 1254 -359 1538 -325
rect 1572 -359 1614 -325
rect 1184 -397 1614 -359
rect 1184 -431 1220 -397
rect 1254 -431 1538 -397
rect 1572 -431 1614 -397
rect 1184 -469 1614 -431
rect 1184 -503 1220 -469
rect 1254 -503 1538 -469
rect 1572 -503 1614 -469
rect 1184 -541 1614 -503
rect 1184 -575 1220 -541
rect 1254 -575 1538 -541
rect 1572 -575 1614 -541
rect 1184 -613 1614 -575
rect 1184 -647 1220 -613
rect 1254 -647 1538 -613
rect 1572 -647 1614 -613
rect 1184 -678 1614 -647
rect 1818 -253 2244 -224
rect 1818 -287 1856 -253
rect 1890 -287 2174 -253
rect 2208 -287 2244 -253
rect 1818 -325 2244 -287
rect 1818 -359 1856 -325
rect 1890 -359 2174 -325
rect 2208 -359 2244 -325
rect 1818 -397 2244 -359
rect 1818 -431 1856 -397
rect 1890 -431 2174 -397
rect 2208 -431 2244 -397
rect 1818 -469 2244 -431
rect 1818 -503 1856 -469
rect 1890 -503 2174 -469
rect 2208 -503 2244 -469
rect 1818 -541 2244 -503
rect 1818 -575 1856 -541
rect 1890 -575 2174 -541
rect 2208 -575 2244 -541
rect 1818 -613 2244 -575
rect 1818 -647 1856 -613
rect 1890 -647 2174 -613
rect 2208 -647 2244 -613
rect 1818 -680 2244 -647
rect -1064 -1089 -940 -1042
rect -1064 -1123 -1024 -1089
rect -990 -1123 -940 -1089
rect -1064 -1161 -940 -1123
rect -1064 -1195 -1024 -1161
rect -990 -1195 -940 -1161
rect -1064 -1233 -940 -1195
rect -1064 -1267 -1024 -1233
rect -990 -1267 -940 -1233
rect -1064 -1305 -940 -1267
rect -1064 -1339 -1024 -1305
rect -990 -1339 -940 -1305
rect -1064 -1377 -940 -1339
rect -1064 -1411 -1024 -1377
rect -990 -1411 -940 -1377
rect -1064 -1449 -940 -1411
rect -1064 -1483 -1024 -1449
rect -990 -1483 -940 -1449
rect -1064 -1676 -940 -1483
rect -766 -1089 -302 -1042
rect -766 -1123 -706 -1089
rect -672 -1123 -388 -1089
rect -354 -1123 -302 -1089
rect -766 -1161 -302 -1123
rect -766 -1195 -706 -1161
rect -672 -1195 -388 -1161
rect -354 -1195 -302 -1161
rect -766 -1233 -302 -1195
rect -766 -1267 -706 -1233
rect -672 -1267 -388 -1233
rect -354 -1267 -302 -1233
rect -766 -1305 -302 -1267
rect -766 -1339 -706 -1305
rect -672 -1339 -388 -1305
rect -354 -1339 -302 -1305
rect -766 -1377 -302 -1339
rect -766 -1411 -706 -1377
rect -672 -1411 -388 -1377
rect -354 -1411 -302 -1377
rect -766 -1449 -302 -1411
rect -766 -1483 -706 -1449
rect -672 -1483 -388 -1449
rect -354 -1483 -302 -1449
rect -766 -1522 -302 -1483
rect -112 -1089 330 -1050
rect -112 -1123 -70 -1089
rect -36 -1123 248 -1089
rect 282 -1123 330 -1089
rect -112 -1161 330 -1123
rect -112 -1195 -70 -1161
rect -36 -1195 248 -1161
rect 282 -1195 330 -1161
rect -112 -1233 330 -1195
rect -112 -1267 -70 -1233
rect -36 -1267 248 -1233
rect 282 -1267 330 -1233
rect -112 -1305 330 -1267
rect -112 -1339 -70 -1305
rect -36 -1339 248 -1305
rect 282 -1339 330 -1305
rect -112 -1377 330 -1339
rect -112 -1411 -70 -1377
rect -36 -1411 248 -1377
rect 282 -1411 330 -1377
rect -112 -1449 330 -1411
rect -112 -1483 -70 -1449
rect -36 -1483 248 -1449
rect 282 -1483 330 -1449
rect -112 -1528 330 -1483
rect 868 -1085 1298 -1046
rect 868 -1119 902 -1085
rect 936 -1119 1220 -1085
rect 1254 -1119 1298 -1085
rect 868 -1157 1298 -1119
rect 868 -1191 902 -1157
rect 936 -1191 1220 -1157
rect 1254 -1191 1298 -1157
rect 868 -1229 1298 -1191
rect 868 -1263 902 -1229
rect 936 -1263 1220 -1229
rect 1254 -1263 1298 -1229
rect 868 -1301 1298 -1263
rect 868 -1335 902 -1301
rect 936 -1335 1220 -1301
rect 1254 -1335 1298 -1301
rect 868 -1373 1298 -1335
rect 868 -1407 902 -1373
rect 936 -1407 1220 -1373
rect 1254 -1407 1298 -1373
rect 868 -1445 1298 -1407
rect 868 -1479 902 -1445
rect 936 -1479 1220 -1445
rect 1254 -1479 1298 -1445
rect 868 -1526 1298 -1479
rect 1504 -1085 1934 -1030
rect 1504 -1119 1538 -1085
rect 1572 -1119 1856 -1085
rect 1890 -1119 1934 -1085
rect 1504 -1157 1934 -1119
rect 1504 -1191 1538 -1157
rect 1572 -1191 1856 -1157
rect 1890 -1191 1934 -1157
rect 1504 -1229 1934 -1191
rect 1504 -1263 1538 -1229
rect 1572 -1263 1856 -1229
rect 1890 -1263 1934 -1229
rect 1504 -1301 1934 -1263
rect 1504 -1335 1538 -1301
rect 1572 -1335 1856 -1301
rect 1890 -1335 1934 -1301
rect 1504 -1373 1934 -1335
rect 1504 -1407 1538 -1373
rect 1572 -1407 1856 -1373
rect 1890 -1407 1934 -1373
rect 1504 -1445 1934 -1407
rect 1504 -1479 1538 -1445
rect 1572 -1479 1856 -1445
rect 1890 -1479 1934 -1445
rect 1504 -1510 1934 -1479
rect 2128 -1085 2256 -1038
rect 2128 -1119 2174 -1085
rect 2208 -1119 2256 -1085
rect 2128 -1157 2256 -1119
rect 2128 -1191 2174 -1157
rect 2208 -1191 2256 -1157
rect 2128 -1229 2256 -1191
rect 2128 -1263 2174 -1229
rect 2208 -1263 2256 -1229
rect 2128 -1301 2256 -1263
rect 2128 -1335 2174 -1301
rect 2208 -1335 2256 -1301
rect 2128 -1373 2256 -1335
rect 2128 -1407 2174 -1373
rect 2208 -1407 2256 -1373
rect 2128 -1445 2256 -1407
rect 2128 -1479 2174 -1445
rect 2208 -1479 2256 -1445
rect -1090 -1708 -940 -1676
rect -744 -1600 -638 -1586
rect -744 -1634 -708 -1600
rect -674 -1634 -638 -1600
rect -1090 -1722 -932 -1708
rect -1090 -1774 -1031 -1722
rect -979 -1774 -932 -1722
rect -1090 -1816 -932 -1774
rect -1072 -2013 -932 -1816
rect -744 -1862 -638 -1634
rect 1830 -1592 1914 -1568
rect 1830 -1626 1850 -1592
rect 1884 -1626 1914 -1592
rect 1830 -1810 1914 -1626
rect 2128 -1679 2256 -1479
rect 2128 -1731 2170 -1679
rect 2222 -1731 2256 -1679
rect 2128 -1734 2256 -1731
rect 1830 -1844 1848 -1810
rect 1882 -1844 1914 -1810
rect 1830 -1862 1914 -1844
rect -744 -1896 -712 -1862
rect -678 -1896 -638 -1862
rect -744 -1908 -638 -1896
rect 1418 -1920 1550 -1918
rect 1322 -1959 1962 -1920
rect -1072 -2047 -1012 -2013
rect -978 -2047 -932 -2013
rect -1072 -2085 -932 -2047
rect -1072 -2119 -1012 -2085
rect -978 -2119 -932 -2085
rect -1072 -2157 -932 -2119
rect -1072 -2191 -1012 -2157
rect -978 -2191 -932 -2157
rect -1072 -2229 -932 -2191
rect -1072 -2263 -1012 -2229
rect -978 -2263 -932 -2229
rect -1072 -2301 -932 -2263
rect -1072 -2335 -1012 -2301
rect -978 -2335 -932 -2301
rect -1072 -2373 -932 -2335
rect -1072 -2407 -1012 -2373
rect -978 -2407 -932 -2373
rect -1072 -2532 -932 -2407
rect -750 -2013 -108 -1974
rect -750 -2047 -694 -2013
rect -660 -2047 -108 -2013
rect -750 -2085 -108 -2047
rect -750 -2119 -694 -2085
rect -660 -2119 -108 -2085
rect -750 -2157 -108 -2119
rect -750 -2191 -694 -2157
rect -660 -2191 -108 -2157
rect -750 -2229 -108 -2191
rect -750 -2263 -694 -2229
rect -660 -2263 -108 -2229
rect -750 -2301 -108 -2263
rect -750 -2335 -694 -2301
rect -660 -2335 -108 -2301
rect -750 -2373 -108 -2335
rect -750 -2407 -694 -2373
rect -660 -2407 -108 -2373
rect -750 -2446 -108 -2407
rect -248 -2604 -108 -2446
rect 1322 -1993 1852 -1959
rect 1886 -1993 1962 -1959
rect 1322 -2031 1962 -1993
rect 1322 -2065 1852 -2031
rect 1886 -2065 1962 -2031
rect 1322 -2103 1962 -2065
rect 1322 -2137 1852 -2103
rect 1886 -2137 1962 -2103
rect 1322 -2175 1962 -2137
rect 1322 -2209 1852 -2175
rect 1886 -2209 1962 -2175
rect 1322 -2247 1962 -2209
rect 1322 -2281 1852 -2247
rect 1886 -2281 1962 -2247
rect 1322 -2319 1962 -2281
rect 1322 -2353 1852 -2319
rect 1886 -2353 1962 -2319
rect 1322 -2392 1962 -2353
rect 2120 -1959 2272 -1734
rect 2120 -1993 2170 -1959
rect 2204 -1993 2272 -1959
rect 2120 -2031 2272 -1993
rect 2120 -2065 2170 -2031
rect 2204 -2065 2272 -2031
rect 2120 -2103 2272 -2065
rect 2120 -2137 2170 -2103
rect 2204 -2137 2272 -2103
rect 2120 -2175 2272 -2137
rect 2120 -2209 2170 -2175
rect 2204 -2209 2272 -2175
rect 2120 -2247 2272 -2209
rect 2120 -2281 2170 -2247
rect 2204 -2281 2272 -2247
rect 2120 -2319 2272 -2281
rect 2120 -2353 2170 -2319
rect 2204 -2353 2272 -2319
rect 1322 -2562 1462 -2392
rect 2120 -2398 2272 -2353
rect -248 -2638 -232 -2604
rect -198 -2638 -160 -2604
rect -126 -2638 -108 -2604
rect -248 -2646 -108 -2638
rect -78 -2606 1288 -2586
rect 1322 -2596 1336 -2562
rect 1370 -2596 1408 -2562
rect 1442 -2596 1462 -2562
rect 1322 -2606 1462 -2596
rect -78 -2618 1248 -2606
rect -78 -2648 173 -2618
rect -78 -2682 -72 -2648
rect -38 -2670 173 -2648
rect 225 -2640 1248 -2618
rect 1282 -2640 1288 -2606
rect 225 -2670 1288 -2640
rect -38 -2682 1288 -2670
rect -248 -2692 -110 -2684
rect -248 -2726 -232 -2692
rect -198 -2726 -160 -2692
rect -126 -2726 -110 -2692
rect -78 -2704 1288 -2682
rect 1324 -2650 1456 -2640
rect 1324 -2684 1336 -2650
rect 1370 -2684 1408 -2650
rect 1442 -2684 1456 -2650
rect -248 -2752 -110 -2726
rect 1324 -2752 1456 -2684
rect -584 -2765 1750 -2752
rect -584 -2770 1258 -2765
rect -584 -2771 130 -2770
rect -584 -2800 -547 -2771
rect -513 -2800 130 -2771
rect -584 -2852 -549 -2800
rect -497 -2805 130 -2800
rect -497 -2839 -310 -2805
rect -276 -2807 -82 -2805
rect -276 -2839 -194 -2807
rect -497 -2841 -194 -2839
rect -160 -2839 -82 -2807
rect -48 -2839 130 -2805
rect -160 -2841 130 -2839
rect -497 -2852 130 -2841
rect -584 -2861 130 -2852
rect -584 -2895 -545 -2861
rect -511 -2884 130 -2861
rect 496 -2773 1258 -2770
rect 496 -2884 696 -2773
rect -511 -2887 696 -2884
rect 1062 -2799 1258 -2773
rect 1292 -2799 1382 -2765
rect 1416 -2799 1486 -2765
rect 1520 -2789 1750 -2765
rect 1520 -2799 1703 -2789
rect 1062 -2823 1703 -2799
rect 1737 -2823 1750 -2789
rect 1062 -2863 1750 -2823
rect 1062 -2887 1703 -2863
rect -511 -2895 1703 -2887
rect -584 -2897 1703 -2895
rect 1737 -2897 1750 -2863
rect -584 -2918 1750 -2897
rect 1802 -4591 2264 -4550
rect -1076 -4645 -614 -4604
rect -1076 -4679 -1012 -4645
rect -978 -4679 -694 -4645
rect -660 -4679 -614 -4645
rect -1076 -4717 -614 -4679
rect -1076 -4751 -1012 -4717
rect -978 -4751 -694 -4717
rect -660 -4751 -614 -4717
rect -1076 -4789 -614 -4751
rect -1076 -4823 -1012 -4789
rect -978 -4823 -694 -4789
rect -660 -4823 -614 -4789
rect -1076 -4861 -614 -4823
rect -1076 -4895 -1012 -4861
rect -978 -4895 -694 -4861
rect -660 -4895 -614 -4861
rect -1076 -4933 -614 -4895
rect -1076 -4967 -1012 -4933
rect -978 -4967 -694 -4933
rect -660 -4967 -614 -4933
rect -1076 -5005 -614 -4967
rect -1076 -5039 -1012 -5005
rect -978 -5039 -694 -5005
rect -660 -5039 -614 -5005
rect 1802 -4625 1852 -4591
rect 1886 -4625 2170 -4591
rect 2204 -4625 2264 -4591
rect 1802 -4663 2264 -4625
rect 1802 -4697 1852 -4663
rect 1886 -4697 2170 -4663
rect 2204 -4697 2264 -4663
rect 1802 -4735 2264 -4697
rect 1802 -4769 1852 -4735
rect 1886 -4769 2170 -4735
rect 2204 -4769 2264 -4735
rect 1802 -4807 2264 -4769
rect 1802 -4841 1852 -4807
rect 1886 -4841 2170 -4807
rect 2204 -4841 2264 -4807
rect 1802 -4879 2264 -4841
rect 1802 -4913 1852 -4879
rect 1886 -4913 2170 -4879
rect 2204 -4913 2264 -4879
rect 1802 -4951 2264 -4913
rect 1802 -4985 1852 -4951
rect 1886 -4985 2170 -4951
rect 2204 -4985 2264 -4951
rect 1802 -5022 2264 -4985
rect -1076 -5076 -614 -5039
<< via1 >>
rect -1224 224 -893 319
rect -903 21 -688 90
rect -624 31 -572 83
rect -1031 -1774 -979 -1722
rect 2170 -1731 2222 -1679
rect 173 -2670 225 -2618
rect -549 -2805 -547 -2800
rect -547 -2805 -513 -2800
rect -513 -2805 -497 -2800
rect -549 -2852 -497 -2805
rect 130 -2884 496 -2770
rect 696 -2887 1062 -2773
<< metal2 >>
rect -1224 319 -893 329
rect -1224 214 -893 224
rect -1364 90 -568 106
rect -1364 21 -903 90
rect -688 83 -568 90
rect -688 31 -624 83
rect -572 31 -568 83
rect -688 21 -568 31
rect -1364 0 -568 21
rect -1364 -120 -1246 0
rect -1364 -2760 -1248 -120
rect 2118 -1677 2284 -1636
rect -1096 -1680 -918 -1678
rect -1096 -1715 -916 -1680
rect -1096 -1722 -1026 -1715
rect -1096 -1774 -1031 -1722
rect -970 -1771 -916 -1715
rect -979 -1774 -916 -1771
rect -1096 -1804 -916 -1774
rect 2118 -1733 2168 -1677
rect 2224 -1733 2284 -1677
rect 2118 -1792 2284 -1733
rect -1096 -1810 -918 -1804
rect 134 -2616 268 -2586
rect 134 -2672 171 -2616
rect 227 -2672 268 -2616
rect 134 -2706 268 -2672
rect -1364 -2770 1082 -2760
rect -1364 -2800 130 -2770
rect -1364 -2852 -549 -2800
rect -497 -2852 130 -2800
rect -1364 -2884 130 -2852
rect 496 -2773 1082 -2770
rect 496 -2884 696 -2773
rect -1364 -2887 696 -2884
rect 1062 -2887 1082 -2773
rect -1364 -2898 1082 -2887
rect -1364 -2900 -1248 -2898
<< via2 >>
rect -1224 224 -893 319
rect -1026 -1722 -970 -1715
rect -1026 -1771 -979 -1722
rect -979 -1771 -970 -1722
rect 2168 -1679 2224 -1677
rect 2168 -1731 2170 -1679
rect 2170 -1731 2222 -1679
rect 2222 -1731 2224 -1679
rect 2168 -1733 2224 -1731
rect 171 -2618 227 -2616
rect 171 -2670 173 -2618
rect 173 -2670 225 -2618
rect 225 -2670 227 -2618
rect 171 -2672 227 -2670
<< metal3 >>
rect -1511 319 -863 339
rect -1511 224 -1224 319
rect -893 224 -863 319
rect -1511 195 -863 224
rect -1318 -2586 -1246 195
rect 2132 -1673 2264 -1636
rect -1088 -1715 -914 -1678
rect -1088 -1779 -1034 -1715
rect -970 -1779 -914 -1715
rect -1088 -1810 -914 -1779
rect 2132 -1737 2161 -1673
rect 2225 -1737 2264 -1673
rect 2132 -1800 2264 -1737
rect -1318 -2616 256 -2586
rect -1318 -2672 171 -2616
rect 227 -2672 256 -2616
rect -1318 -2706 256 -2672
<< via3 >>
rect -1034 -1771 -1026 -1715
rect -1026 -1771 -970 -1715
rect -1034 -1779 -970 -1771
rect 2161 -1677 2225 -1673
rect 2161 -1733 2168 -1677
rect 2168 -1733 2224 -1677
rect 2224 -1733 2225 -1677
rect 2161 -1737 2225 -1733
<< metal4 >>
rect -3498 -1594 -2870 -1384
rect 742 -1673 2278 -1638
rect -1570 -1715 -922 -1676
rect -1570 -1779 -1034 -1715
rect -970 -1779 -922 -1715
rect -1570 -1810 -922 -1779
rect 742 -1737 2161 -1673
rect 2225 -1737 2278 -1673
rect 742 -1796 2278 -1737
rect 742 -2169 880 -1796
rect 742 -2224 879 -2169
rect -1506 -2358 879 -2224
rect -3292 -3018 -2664 -2808
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_0
timestamp 1699818132
transform 1 0 -2274 0 1 -2708
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_1
timestamp 1699818132
transform 1 0 -2284 0 1 -1186
box -786 -640 786 640
use sky130_fd_pr__nfet_01v8_N92D86  sky130_fd_pr__nfet_01v8_N92D86_0
timestamp 1699818132
transform 0 1 -179 -1 0 -2665
box -175 -239 175 239
use sky130_fd_pr__nfet_01v8_N92D86  sky130_fd_pr__nfet_01v8_N92D86_1
timestamp 1699818132
transform 0 1 1389 -1 0 -2623
box -175 -239 175 239
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_0
timestamp 1699818132
transform 0 1 252 -1 0 182
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_1
timestamp 1699818132
transform 0 1 889 -1 0 183
box -211 -319 211 319
use sky130_fd_pr__res_xhigh_po_0p35_RF56VW  sky130_fd_pr__res_xhigh_po_0p35_RF56VW_0
timestamp 1699818132
transform 1 0 -836 0 1 -3526
box -324 -1662 324 1662
use sky130_fd_pr__res_xhigh_po_0p35_RF56VW  sky130_fd_pr__res_xhigh_po_0p35_RF56VW_1
timestamp 1699818132
transform 1 0 2028 0 1 -3472
box -324 -1662 324 1662
use sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ  sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ_0
timestamp 1699818132
transform 1 0 -371 0 1 -870
box -801 -762 801 762
use sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ  sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ_1
timestamp 1699818132
transform 1 0 1555 0 1 -866
box -801 -762 801 762
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699818132
transform 1 0 -634 0 1 56
box -38 -48 314 592
<< labels >>
rlabel metal1 s 71 165 105 199 4 inv_out
rlabel metal1 s 556 342 590 376 4 Vdd
port 1 nsew
rlabel metal1 s -1042 -1798 -962 -1690 4 VP
port 2 nsew
rlabel metal1 s 2154 -1760 2234 -1652 4 VN
port 3 nsew
rlabel metal1 s 532 -2660 590 -2606 4 C1
port 4 nsew
rlabel metal1 s 540 -2860 598 -2806 4 Gnd
port 5 nsew
rlabel metal4 s -3414 -1566 -3306 -1426 4 INP
port 6 nsew
rlabel metal4 s -3180 -2974 -3072 -2834 4 INN
port 7 nsew
<< end >>
