magic
tech sky130A
magscale 1 2
timestamp 1699818132
<< pwell >>
rect -360 640 360 674
rect -360 -640 -326 640
rect 326 -640 360 640
rect -360 -674 360 -640
<< nmoslvt >>
rect -200 -500 200 500
<< ndiff >>
rect -258 459 -200 500
rect -258 425 -246 459
rect -212 425 -200 459
rect -258 391 -200 425
rect -258 357 -246 391
rect -212 357 -200 391
rect -258 323 -200 357
rect -258 289 -246 323
rect -212 289 -200 323
rect -258 255 -200 289
rect -258 221 -246 255
rect -212 221 -200 255
rect -258 187 -200 221
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -221 -200 -187
rect -258 -255 -246 -221
rect -212 -255 -200 -221
rect -258 -289 -200 -255
rect -258 -323 -246 -289
rect -212 -323 -200 -289
rect -258 -357 -200 -323
rect -258 -391 -246 -357
rect -212 -391 -200 -357
rect -258 -425 -200 -391
rect -258 -459 -246 -425
rect -212 -459 -200 -425
rect -258 -500 -200 -459
rect 200 459 258 500
rect 200 425 212 459
rect 246 425 258 459
rect 200 391 258 425
rect 200 357 212 391
rect 246 357 258 391
rect 200 323 258 357
rect 200 289 212 323
rect 246 289 258 323
rect 200 255 258 289
rect 200 221 212 255
rect 246 221 258 255
rect 200 187 258 221
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -221 258 -187
rect 200 -255 212 -221
rect 246 -255 258 -221
rect 200 -289 258 -255
rect 200 -323 212 -289
rect 246 -323 258 -289
rect 200 -357 258 -323
rect 200 -391 212 -357
rect 246 -391 258 -357
rect 200 -425 258 -391
rect 200 -459 212 -425
rect 246 -459 258 -425
rect 200 -500 258 -459
<< ndiffc >>
rect -246 425 -212 459
rect -246 357 -212 391
rect -246 289 -212 323
rect -246 221 -212 255
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect -246 -255 -212 -221
rect -246 -323 -212 -289
rect -246 -391 -212 -357
rect -246 -459 -212 -425
rect 212 425 246 459
rect 212 357 246 391
rect 212 289 246 323
rect 212 221 246 255
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
rect 212 -255 246 -221
rect 212 -323 246 -289
rect 212 -391 246 -357
rect 212 -459 246 -425
<< psubdiff >>
rect -360 640 -255 674
rect -221 640 -187 674
rect -153 640 -119 674
rect -85 640 -51 674
rect -17 640 17 674
rect 51 640 85 674
rect 119 640 153 674
rect 187 640 221 674
rect 255 640 360 674
rect -360 561 -326 640
rect -360 493 -326 527
rect 326 561 360 640
rect -360 425 -326 459
rect -360 357 -326 391
rect -360 289 -326 323
rect -360 221 -326 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -255 -326 -221
rect -360 -323 -326 -289
rect -360 -391 -326 -357
rect -360 -459 -326 -425
rect -360 -527 -326 -493
rect 326 493 360 527
rect 326 425 360 459
rect 326 357 360 391
rect 326 289 360 323
rect 326 221 360 255
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect 326 -255 360 -221
rect 326 -323 360 -289
rect 326 -391 360 -357
rect 326 -459 360 -425
rect -360 -640 -326 -561
rect 326 -527 360 -493
rect 326 -640 360 -561
rect -360 -674 -255 -640
rect -221 -674 -187 -640
rect -153 -674 -119 -640
rect -85 -674 -51 -640
rect -17 -674 17 -640
rect 51 -674 85 -640
rect 119 -674 153 -640
rect 187 -674 221 -640
rect 255 -674 360 -640
<< psubdiffcont >>
rect -255 640 -221 674
rect -187 640 -153 674
rect -119 640 -85 674
rect -51 640 -17 674
rect 17 640 51 674
rect 85 640 119 674
rect 153 640 187 674
rect 221 640 255 674
rect -360 527 -326 561
rect 326 527 360 561
rect -360 459 -326 493
rect -360 391 -326 425
rect -360 323 -326 357
rect -360 255 -326 289
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -360 -289 -326 -255
rect -360 -357 -326 -323
rect -360 -425 -326 -391
rect -360 -493 -326 -459
rect 326 459 360 493
rect 326 391 360 425
rect 326 323 360 357
rect 326 255 360 289
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect 326 -289 360 -255
rect 326 -357 360 -323
rect 326 -425 360 -391
rect 326 -493 360 -459
rect -360 -561 -326 -527
rect 326 -561 360 -527
rect -255 -674 -221 -640
rect -187 -674 -153 -640
rect -119 -674 -85 -640
rect -51 -674 -17 -640
rect 17 -674 51 -640
rect 85 -674 119 -640
rect 153 -674 187 -640
rect 221 -674 255 -640
<< poly >>
rect -200 572 200 588
rect -200 538 -153 572
rect -119 538 -85 572
rect -51 538 -17 572
rect 17 538 51 572
rect 85 538 119 572
rect 153 538 200 572
rect -200 500 200 538
rect -200 -538 200 -500
rect -200 -572 -153 -538
rect -119 -572 -85 -538
rect -51 -572 -17 -538
rect 17 -572 51 -538
rect 85 -572 119 -538
rect 153 -572 200 -538
rect -200 -588 200 -572
<< polycont >>
rect -153 538 -119 572
rect -85 538 -51 572
rect -17 538 17 572
rect 51 538 85 572
rect 119 538 153 572
rect -153 -572 -119 -538
rect -85 -572 -51 -538
rect -17 -572 17 -538
rect 51 -572 85 -538
rect 119 -572 153 -538
<< locali >>
rect -360 640 -255 674
rect -221 640 -187 674
rect -153 640 -119 674
rect -85 640 -51 674
rect -17 640 17 674
rect 51 640 85 674
rect 119 640 153 674
rect 187 640 221 674
rect 255 640 360 674
rect -360 561 -326 640
rect -200 538 -153 572
rect -119 538 -85 572
rect -51 538 -17 572
rect 17 538 51 572
rect 85 538 119 572
rect 153 538 200 572
rect 326 561 360 640
rect -360 493 -326 527
rect -360 425 -326 459
rect -360 357 -326 391
rect -360 289 -326 323
rect -360 221 -326 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -255 -326 -221
rect -360 -323 -326 -289
rect -360 -391 -326 -357
rect -360 -459 -326 -425
rect -360 -527 -326 -493
rect -246 459 -212 504
rect -246 391 -212 425
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect -246 -425 -212 -391
rect -246 -504 -212 -459
rect 212 459 246 504
rect 212 391 246 425
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
rect 212 -425 246 -391
rect 212 -504 246 -459
rect 326 493 360 527
rect 326 425 360 459
rect 326 357 360 391
rect 326 289 360 323
rect 326 221 360 255
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect 326 -255 360 -221
rect 326 -323 360 -289
rect 326 -391 360 -357
rect 326 -459 360 -425
rect 326 -527 360 -493
rect -360 -640 -326 -561
rect -200 -572 -153 -538
rect -119 -572 -85 -538
rect -51 -572 -17 -538
rect 17 -572 51 -538
rect 85 -572 119 -538
rect 153 -572 200 -538
rect 326 -640 360 -561
rect -360 -674 -255 -640
rect -221 -674 -187 -640
rect -153 -674 -119 -640
rect -85 -674 -51 -640
rect -17 -674 17 -640
rect 51 -674 85 -640
rect 119 -674 153 -640
rect 187 -674 221 -640
rect 255 -674 360 -640
<< properties >>
string FIXED_BBOX -342 -656 342 656
<< end >>
